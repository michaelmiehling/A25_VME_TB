-- megafunction wizard: %ALTASMI_PARALLEL%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTASMI_PARALLEL 

-- ============================================================
-- File Name: z126_01_pasmi_sim_m25p32_2.vhd
-- Megafunction Name(s):
-- 			ALTASMI_PARALLEL
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 11.1 Build 259 01/25/2012 SP 2 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2011 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altasmi_parallel CBX_AUTO_BLACKBOX="ALL" DATA_WIDTH="STANDARD" DEVICE_FAMILY="Cyclone III" EPCS_TYPE="EPCS16" PAGE_SIZE=256 PORT_BULK_ERASE="PORT_USED" PORT_EN4B_ADDR="PORT_UNUSED" PORT_FAST_READ="PORT_USED" PORT_ILLEGAL_ERASE="PORT_USED" PORT_ILLEGAL_WRITE="PORT_USED" PORT_RDID_OUT="PORT_USED" PORT_READ_ADDRESS="PORT_UNUSED" PORT_READ_RDID="PORT_USED" PORT_READ_SID="PORT_UNUSED" PORT_READ_STATUS="PORT_USED" PORT_SECTOR_ERASE="PORT_USED" PORT_SECTOR_PROTECT="PORT_USED" PORT_SHIFT_BYTES="PORT_USED" PORT_WREN="PORT_USED" PORT_WRITE="PORT_USED" USE_EAB="ON" addr bulk_erase busy clkin data_valid datain dataout fast_read illegal_erase illegal_write rden rdid_out read_rdid read_status sector_erase sector_protect shift_bytes status_out wren write INTENDED_DEVICE_FAMILY="Cyclone III" ALTERA_INTERNAL_OPTIONS=SUPPRESS_DA_RULE_INTERNAL=C106
--VERSION_BEGIN 11.1SP2 cbx_a_gray2bin 2012:01:25:21:14:55:SJ cbx_a_graycounter 2012:01:25:21:14:55:SJ cbx_altasmi_parallel 2012:01:25:21:14:55:SJ cbx_altdpram 2012:01:25:21:14:55:SJ cbx_altsyncram 2012:01:25:21:14:56:SJ cbx_cyclone 2012:01:25:21:14:56:SJ cbx_cycloneii 2012:01:25:21:14:56:SJ cbx_fifo_common 2012:01:25:21:14:55:SJ cbx_lpm_add_sub 2012:01:25:21:14:56:SJ cbx_lpm_compare 2012:01:25:21:14:56:SJ cbx_lpm_counter 2012:01:25:21:14:56:SJ cbx_lpm_decode 2012:01:25:21:14:56:SJ cbx_lpm_mux 2012:01:25:21:14:56:SJ cbx_mgl 2012:01:25:21:17:49:SJ cbx_scfifo 2012:01:25:21:14:56:SJ cbx_stratix 2012:01:25:21:14:56:SJ cbx_stratixii 2012:01:25:21:14:56:SJ cbx_stratixiii 2012:01:25:21:14:56:SJ cbx_stratixv 2012:01:25:21:14:56:SJ cbx_util_mgl 2012:01:25:21:14:56:SJ  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY cycloneii;
 USE cycloneii.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = a_graycounter 5 cycloneii_asmiblock 1 lpm_compare 2 lpm_counter 2 lut 70 mux21 2 reg 147 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  z126_01_pasmi_sim_m25p32_altasmi_parallel_l2q2 IS 
	 PORT 
	 ( 
		 addr	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 bulk_erase	:	IN  STD_LOGIC := '0';
		 busy	:	OUT  STD_LOGIC;
		 clkin	:	IN  STD_LOGIC;
		 data_valid	:	OUT  STD_LOGIC;
		 datain	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 dataout	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 fast_read	:	IN  STD_LOGIC := '0';
		 illegal_erase	:	OUT  STD_LOGIC;
		 illegal_write	:	OUT  STD_LOGIC;
		 rden	:	IN  STD_LOGIC;
		 rdid_out	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 read_rdid	:	IN  STD_LOGIC := '0';
		 read_status	:	IN  STD_LOGIC := '0';
		 sector_erase	:	IN  STD_LOGIC := '0';
		 sector_protect	:	IN  STD_LOGIC := '0';
		 shift_bytes	:	IN  STD_LOGIC := '0';
		 status_out	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 wren	:	IN  STD_LOGIC := '1';
		 write	:	IN  STD_LOGIC := '0'
	 ); 
 END z126_01_pasmi_sim_m25p32_altasmi_parallel_l2q2;

 ARCHITECTURE RTL OF z126_01_pasmi_sim_m25p32_altasmi_parallel_l2q2 IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "SUPPRESS_DA_RULE_INTERNAL=C106";

	 SIGNAL  wire_addbyte_cntr_w_lg_w_q_range137w142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_lg_w_q_range140w141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w135w136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_clock	:	STD_LOGIC;
	 SIGNAL  wire_addbyte_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_q_range140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_q_range137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_lg_w_q_range99w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_lg_w_q_range97w98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_in_operation44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_q_range97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_q_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_spstage_cntr_w_lg_w_q_range598w599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_spstage_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_do_sec_prot595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_spstage_cntr_clock	:	STD_LOGIC;
	 SIGNAL  wire_spstage_cntr_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_spstage_cntr_w_q_range596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_spstage_cntr_w_q_range598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w247w248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w92w244w245w246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w92w249w250w251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w90w91w257w258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w94w322w323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w269w270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w244w245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w249w250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w90w91w257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range89w94w322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range89w92w269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range89w92w244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range89w92w249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range89w92w135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w93w107w108w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range88w93w107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range89w90w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range89w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range89w92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w93w107w108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range88w93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range89w90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w82w83w84w85w86w87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_q_range88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_q_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_lg_w_q_range494w495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_lg_w_q_range492w493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w490w491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_clock	:	STD_LOGIC;
	 SIGNAL  wire_wrstage_cntr_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_q_range492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_q_range494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cycloneii_asmiblock3_data0out	:	STD_LOGIC;
	 SIGNAL	 add_msb_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_add_msb_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_addr_reg_d	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL	 addr_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_addr_reg_ena	:	STD_LOGIC_VECTOR(23 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w535w536w537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w535w536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range512w518w524w525w526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range512w518w524w529w530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range512w518w524w529w534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_lg_w_q_range512w513w514w515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_lg_w_q_range512w518w524w525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_lg_w_q_range512w518w524w529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_q_range512w513w514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_q_range512w518w519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_q_range512w518w524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_q_range512w513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_q_range512w518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range301w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL	 wire_asmi_opcode_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 asmi_opcode_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_asmi_opcode_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_asmi_opcode_reg_w_q_range147w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL	 buf_empty_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 bulk_erase_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_bulk_erase_reg_ena	:	STD_LOGIC;
	 SIGNAL	 busy_delay_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 busy_det_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_addmsb_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_endrbyte_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_clr_endrbyte_reg_w_lg_q388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 clr_rdid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_rdid_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_read_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_rstat_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_rstat_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_secprot_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_secprot_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_write_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_write_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cnt_bfend_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 do_wrmemadd_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dvalid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dvalid_reg_ena	:	STD_LOGIC;
	 SIGNAL	 dvalid_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end1_cyc_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end1_cyc_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_op_hdlyreg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_op_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_opfdly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_pgwrop_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_end_pgwrop_reg_ena	:	STD_LOGIC;
	 SIGNAL	 end_rbyte_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_end_rbyte_reg_ena	:	STD_LOGIC;
	 SIGNAL	 end_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 fast_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_fast_read_reg_ena	:	STD_LOGIC;
	 SIGNAL	 ill_erase_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 ill_write_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 illegal_erase_dly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 illegal_write_dly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 max_cnt_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 maxcnt_shift_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 maxcnt_shift_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 ncs_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_ncs_reg_ena	:	STD_LOGIC;
	 SIGNAL  wire_ncs_reg_w_lg_q291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_pgwrbuf_dataout_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 pgwrbuf_dataout	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_pgwrbuf_dataout_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_pgwrbuf_dataout_w_q_range438w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL	 power_up_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rdid_out_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_bufdly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_data_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 read_data_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_data_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 wire_read_dout_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 read_dout_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_dout_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 read_rdid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_status_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sec_erase_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_sec_erase_reg_ena	:	STD_LOGIC;
	 SIGNAL	 sec_prot_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_sec_prot_reg_ena	:	STD_LOGIC;
	 SIGNAL	 shftpgwr_data_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 shift_op_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sprot_rstat_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage2_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage3_dly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage3_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage4_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 start_sppoll_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_start_sppoll_reg_ena	:	STD_LOGIC;
	 SIGNAL	 start_sppoll_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 start_wrpoll_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_start_wrpoll_reg_ena	:	STD_LOGIC;
	 SIGNAL	 start_wrpoll_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_statreg_int_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 statreg_int	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_statreg_int_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 wire_statreg_out_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 statreg_out	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_statreg_out_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 streg_datain_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_streg_datain_reg_ena	:	STD_LOGIC;
	 SIGNAL	 write_prot_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_write_prot_reg_ena	:	STD_LOGIC;
	 SIGNAL	 write_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_write_reg_ena	:	STD_LOGIC;
	 SIGNAL	 write_rstat_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_wrstat_dreg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 wrstat_dreg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_wrstat_dreg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_wrstat_dreg_w_q_range602w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_cmpr5_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr5_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_cmpr5_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_cmpr6_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr6_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_cmpr6_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_shift_bytes_wire434w450w451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_q	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_read_cntr_q	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL	wire_mux211_dataout	:	STD_LOGIC;
	 SIGNAL	wire_mux212_dataout	:	STD_LOGIC;
	 SIGNAL  wire_scfifo4_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_scfifo4_q	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_scfifo4_rdreq	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_read_buf436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_scfifo4_wrreq	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_shift_bytes_wire434w435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_scfifo4_w_q_range441w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_scfifo4_w_q_range446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w413w414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_end_operation409w410w411w412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode158w159w160w210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode158w159w160w161w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode163w164w165w212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode163w164w165w166w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode182w183w184w222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode182w183w184w185w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read274w275w276w277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write408w581w582w583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w586w587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read330w374w375w376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_sec_erase318w319w320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_sec_prot612w613w614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_end_operation409w410w411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode158w159w160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode163w164w165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode182w183w184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read274w275w276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read274w275w321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write408w581w582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read330w374w375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_4baddr150w151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_polling420w421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_sec_erase318w319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_sec_prot612w613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write171w172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write56w253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_end_operation409w410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode152w206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode152w153w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode173w216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode173w174w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode158w159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode176w218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode176w177w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode179w220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode179w180w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode187w224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode187w188w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode190w226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode190w191w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode168w214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode168w169w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode163w164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode182w183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode155w208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode155w156w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_reach_max_cnt484w485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_start_poll259w260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read274w275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write408w581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_bufdly439w440w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write65w66w499w585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write65w66w488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write65w66w67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read330w374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write65w311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_end_operation422w423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rden_wire315w316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_4baddr150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_bulk_erase254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_polling420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_erase318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_prot600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_prot612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_prot621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_operation409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy304w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy605w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_reach_max_cnt484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly442w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_opcode148w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire302w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire603w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_start_poll259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_wren_wire615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write56w272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp0_wire516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp1_wire511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp2_wire522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_buf_empty553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_busy_wire2w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clkin_wire42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_4baddr404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_bulk_erase406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_fast_read273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_memadd327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_polling268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_rdid45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_erase407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_prot405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_wren47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_add_cycle75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_fast_read69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_ophdly43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_pgwr_data55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_read72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rden_wire389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reach_max_cnt449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_rdid_wire11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_sid_wire10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_status_wire26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sec_erase_wire29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sec_protect_wire14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_st_busy_wire102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_prot_true487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_wire21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range61w62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w586w587w588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode190w226w227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode190w191w192w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write65w66w488w489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write65w311w312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_rden_wire315w316w317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_not_busy304w305w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_not_busy605w606w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_bufdly442w443w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage4_wire343w344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_wren_wire615w616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode190w226w227w228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode190w191w192w193w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write65w311w312w313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w194w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w229w230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w194w195w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w229w230w231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w194w195w196w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w229w230w231w232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w194w195w196w197w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w229w230w231w232w233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w194w195w196w197w198w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w229w230w231w232w233w234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w194w195w196w197w198w199w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w200w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w235w236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w200w201w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w200w201w202w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read_sid130w131w132w133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read330w331w332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_sid130w131w132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write65w66w499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read330w342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read330w331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_sid130w131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_sec_erase501w502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write65w66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_data0out_wire346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_4baddr255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_sid130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_erase501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_wren256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_operation422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rden_wire315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range453w456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range457w459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range460w462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range463w465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range466w468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range469w471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range472w474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range475w477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  b4addr_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  be_write_prot :	STD_LOGIC;
	 SIGNAL  berase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  bp0_wire :	STD_LOGIC;
	 SIGNAL  bp1_wire :	STD_LOGIC;
	 SIGNAL  bp2_wire :	STD_LOGIC;
	 SIGNAL  bp3_wire :	STD_LOGIC;
	 SIGNAL  buf_empty :	STD_LOGIC;
	 SIGNAL  bulk_erase_wire :	STD_LOGIC;
	 SIGNAL  busy_wire :	STD_LOGIC;
	 SIGNAL  clkin_wire :	STD_LOGIC;
	 SIGNAL  clr_rdid_wire :	STD_LOGIC;
	 SIGNAL  clr_read_wire :	STD_LOGIC;
	 SIGNAL  clr_rstat_wire :	STD_LOGIC;
	 SIGNAL  clr_secprot_wire :	STD_LOGIC;
	 SIGNAL  clr_write_wire :	STD_LOGIC;
	 SIGNAL  cnt_bfend_wire_in :	STD_LOGIC;
	 SIGNAL  data0out_wire :	STD_LOGIC;
	 SIGNAL  data_valid_wire :	STD_LOGIC;
	 SIGNAL  dataout_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  do_4baddr :	STD_LOGIC;
	 SIGNAL  do_bulk_erase :	STD_LOGIC;
	 SIGNAL  do_fast_read :	STD_LOGIC;
	 SIGNAL  do_memadd :	STD_LOGIC;
	 SIGNAL  do_polling :	STD_LOGIC;
	 SIGNAL  do_read :	STD_LOGIC;
	 SIGNAL  do_read_rdid :	STD_LOGIC;
	 SIGNAL  do_read_sid :	STD_LOGIC;
	 SIGNAL  do_read_stat :	STD_LOGIC;
	 SIGNAL  do_sec_erase :	STD_LOGIC;
	 SIGNAL  do_sec_prot :	STD_LOGIC;
	 SIGNAL  do_secprot_wren :	STD_LOGIC;
	 SIGNAL  do_sprot_polling :	STD_LOGIC;
	 SIGNAL  do_sprot_rstat :	STD_LOGIC;
	 SIGNAL  do_wren :	STD_LOGIC;
	 SIGNAL  do_write :	STD_LOGIC;
	 SIGNAL  do_write_polling :	STD_LOGIC;
	 SIGNAL  do_write_rstat :	STD_LOGIC;
	 SIGNAL  do_write_wren :	STD_LOGIC;
	 SIGNAL  dummy_read_buf :	STD_LOGIC;
	 SIGNAL  end1_cyc_dlyncs_in_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_gen_cntr_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_normal_in_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_reg_in_wire :	STD_LOGIC;
	 SIGNAL  end_add_cycle :	STD_LOGIC;
	 SIGNAL  end_add_cycle_mux_datab_wire :	STD_LOGIC;
	 SIGNAL  end_fast_read :	STD_LOGIC;
	 SIGNAL  end_one_cyc_pos :	STD_LOGIC;
	 SIGNAL  end_one_cycle :	STD_LOGIC;
	 SIGNAL  end_operation :	STD_LOGIC;
	 SIGNAL  end_opfdly :	STD_LOGIC;
	 SIGNAL  end_ophdly :	STD_LOGIC;
	 SIGNAL  end_pgwr_data :	STD_LOGIC;
	 SIGNAL  end_read :	STD_LOGIC;
	 SIGNAL  end_read_byte :	STD_LOGIC;
	 SIGNAL  end_wrstage :	STD_LOGIC;
	 SIGNAL  fast_read_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  fast_read_wire :	STD_LOGIC;
	 SIGNAL  ill_erase_wire :	STD_LOGIC;
	 SIGNAL  ill_write_wire :	STD_LOGIC;
	 SIGNAL  illegal_erase_b4out_wire :	STD_LOGIC;
	 SIGNAL  illegal_write_b4out_wire :	STD_LOGIC;
	 SIGNAL  in_operation :	STD_LOGIC;
	 SIGNAL  load_opcode :	STD_LOGIC;
	 SIGNAL  memadd_sdoin :	STD_LOGIC;
	 SIGNAL  not_busy :	STD_LOGIC;
	 SIGNAL  oe_wire :	STD_LOGIC;
	 SIGNAL  page_size_wire :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  pagewr_buf_not_empty :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  rden_wire :	STD_LOGIC;
	 SIGNAL  rdid_load :	STD_LOGIC;
	 SIGNAL  rdid_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  reach_max_cnt :	STD_LOGIC;
	 SIGNAL  read_buf :	STD_LOGIC;
	 SIGNAL  read_bufdly :	STD_LOGIC;
	 SIGNAL  read_data_reg_in_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_rdid_wire :	STD_LOGIC;
	 SIGNAL  read_sid_wire :	STD_LOGIC;
	 SIGNAL  read_status_wire :	STD_LOGIC;
	 SIGNAL  read_wire :	STD_LOGIC;
	 SIGNAL  rsid_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rsid_sdoin :	STD_LOGIC;
	 SIGNAL  rstat_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  scein_wire :	STD_LOGIC;
	 SIGNAL  sdoin_wire :	STD_LOGIC;
	 SIGNAL  sec_erase_wire :	STD_LOGIC;
	 SIGNAL  sec_protect_wire :	STD_LOGIC;
	 SIGNAL  secprot_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  secprot_sdoin :	STD_LOGIC;
	 SIGNAL  serase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  shift_bytes_wire :	STD_LOGIC;
	 SIGNAL  shift_opcode :	STD_LOGIC;
	 SIGNAL  shift_opdata :	STD_LOGIC;
	 SIGNAL  shift_pgwr_data :	STD_LOGIC;
	 SIGNAL  st_busy_wire :	STD_LOGIC;
	 SIGNAL  stage2_wire :	STD_LOGIC;
	 SIGNAL  stage3_wire :	STD_LOGIC;
	 SIGNAL  stage4_wire :	STD_LOGIC;
	 SIGNAL  start_poll :	STD_LOGIC;
	 SIGNAL  start_sppoll :	STD_LOGIC;
	 SIGNAL  start_wrpoll :	STD_LOGIC;
	 SIGNAL  to_sdoin_wire :	STD_LOGIC;
	 SIGNAL  wren_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wren_wire :	STD_LOGIC;
	 SIGNAL  write_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  write_prot_true :	STD_LOGIC;
	 SIGNAL  write_sdoin :	STD_LOGIC;
	 SIGNAL  write_wire :	STD_LOGIC;
	 SIGNAL  wire_w_addr_range308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_addr_range303w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_b4addr_opcode_range205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_b4addr_opcode_range149w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_berase_opcode_range209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_berase_opcode_range157w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_datain_range609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datain_range604w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_dataout_wire_range345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_fast_read_opcode_range217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_fast_read_opcode_range175w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdid_opcode_range223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdid_opcode_range186w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_read_opcode_range219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_read_opcode_range178w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rsid_opcode_range225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rsid_opcode_range189w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rstat_opcode_range213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rstat_opcode_range167w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_secprot_opcode_range221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_secprot_opcode_range181w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_serase_opcode_range211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_serase_opcode_range162w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_wren_opcode_range207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wren_opcode_range154w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_write_opcode_range215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_write_opcode_range170w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 COMPONENT  a_graycounter
	 GENERIC 
	 (
		PVALUE	:	NATURAL := 0;
		WIDTH	:	NATURAL := 8;
		lpm_type	:	STRING := "a_graycounter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		q	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		qbin	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  cycloneii_asmiblock
	 PORT
	 ( 
		data0out	:	OUT STD_LOGIC;
		dclkin	:	IN STD_LOGIC;
		oe	:	IN STD_LOGIC := '1';
		scein	:	IN STD_LOGIC;
		sdoin	:	IN STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  scfifo
	 GENERIC 
	 (
		ADD_RAM_OUTPUT_REGISTER	:	STRING := "OFF";
		ALLOW_RWCYCLE_WHEN_FULL	:	STRING := "OFF";
		ALMOST_EMPTY_VALUE	:	NATURAL := 0;
		ALMOST_FULL_VALUE	:	NATURAL := 0;
		LPM_NUMWORDS	:	NATURAL;
		LPM_SHOWAHEAD	:	STRING := "OFF";
		LPM_WIDTH	:	NATURAL;
		LPM_WIDTHU	:	NATURAL := 1;
		OVERFLOW_CHECKING	:	STRING := "ON";
		UNDERFLOW_CHECKING	:	STRING := "ON";
		USE_EAB	:	STRING := "ON";
		lpm_type	:	STRING := "scfifo"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		almost_empty	:	OUT STD_LOGIC;
		almost_full	:	OUT STD_LOGIC;
		clock	:	IN STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		empty	:	OUT STD_LOGIC;
		full	:	OUT STD_LOGIC;
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		rdreq	:	IN STD_LOGIC;
		sclr	:	IN STD_LOGIC := '0';
		usedw	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHU-1 DOWNTO 0);
		wrreq	:	IN STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w413w414w(0) <= wire_w413w(0) AND wire_w_lg_do_4baddr404w(0);
	wire_w413w(0) <= wire_w_lg_w_lg_w_lg_w_lg_end_operation409w410w411w412w(0) AND wire_w_lg_do_sec_prot405w(0);
	wire_w584w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write408w581w582w583w(0) AND end_operation;
	wire_w377w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read330w374w375w376w(0) AND end_read_byte;
	wire_w_lg_w_lg_w_lg_w_lg_end_operation409w410w411w412w(0) <= wire_w_lg_w_lg_w_lg_end_operation409w410w411w(0) AND wire_w_lg_do_bulk_erase406w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode158w159w160w210w(0) <= wire_w_lg_w_lg_w_lg_load_opcode158w159w160w(0) AND wire_w_berase_opcode_range209w(0);
	loop0 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode158w159w160w161w(i) <= wire_w_lg_w_lg_w_lg_load_opcode158w159w160w(0) AND wire_w_berase_opcode_range157w(i);
	END GENERATE loop0;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode163w164w165w212w(0) <= wire_w_lg_w_lg_w_lg_load_opcode163w164w165w(0) AND wire_w_serase_opcode_range211w(0);
	loop1 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode163w164w165w166w(i) <= wire_w_lg_w_lg_w_lg_load_opcode163w164w165w(0) AND wire_w_serase_opcode_range162w(i);
	END GENERATE loop1;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode182w183w184w222w(0) <= wire_w_lg_w_lg_w_lg_load_opcode182w183w184w(0) AND wire_w_secprot_opcode_range221w(0);
	loop2 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode182w183w184w185w(i) <= wire_w_lg_w_lg_w_lg_load_opcode182w183w184w(0) AND wire_w_secprot_opcode_range181w(i);
	END GENERATE loop2;
	wire_w_lg_w_lg_w_lg_w_lg_do_read274w275w276w277w(0) <= wire_w_lg_w_lg_w_lg_do_read274w275w276w(0) AND end_one_cycle;
	wire_w_lg_w_lg_w_lg_w_lg_do_write408w581w582w583w(0) <= wire_w_lg_w_lg_w_lg_do_write408w581w582w(0) AND wire_w_lg_do_4baddr404w(0);
	wire_w_lg_w586w587w(0) <= wire_w586w(0) AND end_operation;
	wire_w_lg_w_lg_w_lg_w_lg_do_read330w374w375w376w(0) <= wire_w_lg_w_lg_w_lg_do_read330w374w375w(0) AND end_one_cyc_pos;
	wire_w_lg_w_lg_w_lg_do_sec_erase318w319w320w(0) <= wire_w_lg_w_lg_do_sec_erase318w319w(0) AND end_operation;
	wire_w_lg_w_lg_w_lg_do_sec_prot612w613w614w(0) <= wire_w_lg_w_lg_do_sec_prot612w613w(0) AND wire_spstage_cntr_w_q_range596w(0);
	wire_w_lg_w_lg_w_lg_end_operation409w410w411w(0) <= wire_w_lg_w_lg_end_operation409w410w(0) AND wire_w_lg_do_sec_erase407w(0);
	wire_w_lg_w_lg_w_lg_load_opcode158w159w160w(0) <= wire_w_lg_w_lg_load_opcode158w159w(0) AND wire_w_lg_do_read_stat46w(0);
	wire_w_lg_w_lg_w_lg_load_opcode163w164w165w(0) <= wire_w_lg_w_lg_load_opcode163w164w(0) AND wire_w_lg_do_read_stat46w(0);
	wire_w_lg_w_lg_w_lg_load_opcode182w183w184w(0) <= wire_w_lg_w_lg_load_opcode182w183w(0) AND wire_w_lg_do_read_stat46w(0);
	wire_w_lg_w_lg_w_lg_do_read274w275w276w(0) <= wire_w_lg_w_lg_do_read274w275w(0) AND wire_w_lg_w_lg_do_write56w272w(0);
	wire_w_lg_w_lg_w_lg_do_read274w275w321w(0) <= wire_w_lg_w_lg_do_read274w275w(0) AND clr_write_wire;
	wire_w_lg_w_lg_w_lg_do_write408w581w582w(0) <= wire_w_lg_w_lg_do_write408w581w(0) AND wire_w_lg_do_bulk_erase406w(0);
	wire_w586w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write65w66w499w585w(0) AND wire_wrstage_cntr_w_lg_w_q_range492w493w(0);
	wire_w_lg_w_lg_w_lg_do_read330w374w375w(0) <= wire_w_lg_w_lg_do_read330w374w(0) AND wire_stage_cntr_w_lg_w_q_range88w93w(0);
	wire_w_lg_w_lg_do_4baddr150w151w(0) <= wire_w_lg_do_4baddr150w(0) AND wire_w_lg_do_wren47w(0);
	wire_w_lg_w_lg_do_polling420w421w(0) <= wire_w_lg_do_polling420w(0) AND stage3_dly_reg;
	wire_w_lg_w_lg_do_sec_erase318w319w(0) <= wire_w_lg_do_sec_erase318w(0) AND wire_w_lg_do_read_stat46w(0);
	wire_w_lg_w_lg_do_sec_prot612w613w(0) <= wire_w_lg_do_sec_prot612w(0) AND wire_spstage_cntr_w_lg_w_q_range598w599w(0);
	wire_w_lg_w_lg_do_write171w172w(0) <= wire_w_lg_do_write171w(0) AND wire_w_lg_do_wren47w(0);
	wire_w_lg_w_lg_do_write56w253w(0) <= wire_w_lg_do_write56w(0) AND end_pgwr_data;
	wire_w_lg_w_lg_end_operation409w410w(0) <= wire_w_lg_end_operation409w(0) AND wire_w_lg_do_write408w(0);
	wire_w_lg_w_lg_load_opcode152w206w(0) <= wire_w_lg_load_opcode152w(0) AND wire_w_b4addr_opcode_range205w(0);
	loop3 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode152w153w(i) <= wire_w_lg_load_opcode152w(0) AND wire_w_b4addr_opcode_range149w(i);
	END GENERATE loop3;
	wire_w_lg_w_lg_load_opcode173w216w(0) <= wire_w_lg_load_opcode173w(0) AND wire_w_write_opcode_range215w(0);
	loop4 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode173w174w(i) <= wire_w_lg_load_opcode173w(0) AND wire_w_write_opcode_range170w(i);
	END GENERATE loop4;
	wire_w_lg_w_lg_load_opcode158w159w(0) <= wire_w_lg_load_opcode158w(0) AND wire_w_lg_do_wren47w(0);
	wire_w_lg_w_lg_load_opcode176w218w(0) <= wire_w_lg_load_opcode176w(0) AND wire_w_fast_read_opcode_range217w(0);
	loop5 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode176w177w(i) <= wire_w_lg_load_opcode176w(0) AND wire_w_fast_read_opcode_range175w(i);
	END GENERATE loop5;
	wire_w_lg_w_lg_load_opcode179w220w(0) <= wire_w_lg_load_opcode179w(0) AND wire_w_read_opcode_range219w(0);
	loop6 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode179w180w(i) <= wire_w_lg_load_opcode179w(0) AND wire_w_read_opcode_range178w(i);
	END GENERATE loop6;
	wire_w_lg_w_lg_load_opcode187w224w(0) <= wire_w_lg_load_opcode187w(0) AND wire_w_rdid_opcode_range223w(0);
	loop7 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode187w188w(i) <= wire_w_lg_load_opcode187w(0) AND wire_w_rdid_opcode_range186w(i);
	END GENERATE loop7;
	wire_w_lg_w_lg_load_opcode190w226w(0) <= wire_w_lg_load_opcode190w(0) AND wire_w_rsid_opcode_range225w(0);
	loop8 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode190w191w(i) <= wire_w_lg_load_opcode190w(0) AND wire_w_rsid_opcode_range189w(i);
	END GENERATE loop8;
	wire_w_lg_w_lg_load_opcode168w214w(0) <= wire_w_lg_load_opcode168w(0) AND wire_w_rstat_opcode_range213w(0);
	loop9 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode168w169w(i) <= wire_w_lg_load_opcode168w(0) AND wire_w_rstat_opcode_range167w(i);
	END GENERATE loop9;
	wire_w_lg_w_lg_load_opcode163w164w(0) <= wire_w_lg_load_opcode163w(0) AND wire_w_lg_do_wren47w(0);
	wire_w_lg_w_lg_load_opcode182w183w(0) <= wire_w_lg_load_opcode182w(0) AND wire_w_lg_do_wren47w(0);
	wire_w_lg_w_lg_load_opcode155w208w(0) <= wire_w_lg_load_opcode155w(0) AND wire_w_wren_opcode_range207w(0);
	loop10 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode155w156w(i) <= wire_w_lg_load_opcode155w(0) AND wire_w_wren_opcode_range154w(i);
	END GENERATE loop10;
	wire_w_lg_w_lg_reach_max_cnt484w485w(0) <= wire_w_lg_reach_max_cnt484w(0) AND wren_wire;
	wire_w_lg_w_lg_start_poll259w260w(0) <= wire_w_lg_start_poll259w(0) AND do_polling;
	wire_w_lg_w_lg_do_read274w275w(0) <= wire_w_lg_do_read274w(0) AND wire_w_lg_do_fast_read273w(0);
	wire_w_lg_w_lg_do_write408w581w(0) <= wire_w_lg_do_write408w(0) AND wire_w_lg_do_sec_erase407w(0);
	loop11 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_read_bufdly439w440w(i) <= wire_w_lg_read_bufdly439w(0) AND wire_pgwrbuf_dataout_w_q_range438w(i);
	END GENERATE loop11;
	wire_w490w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write65w66w488w489w(0) AND end_wrstage;
	wire_w_lg_w_lg_w_lg_w_lg_do_write65w66w499w585w(0) <= wire_w_lg_w_lg_w_lg_do_write65w66w499w(0) AND wire_wrstage_cntr_w_q_range494w(0);
	wire_w_lg_w_lg_w_lg_do_write65w66w488w(0) <= wire_w_lg_w_lg_do_write65w66w(0) AND wire_w_lg_write_prot_true487w(0);
	wire_w_lg_w_lg_w_lg_do_write65w66w67w(0) <= wire_w_lg_w_lg_do_write65w66w(0) AND write_prot_true;
	wire_w_lg_w_lg_do_read330w374w(0) <= wire_w_lg_do_read330w(0) AND wire_stage_cntr_w_q_range89w(0);
	wire_w_lg_w_lg_do_write65w311w(0) <= wire_w_lg_do_write65w(0) AND do_memadd;
	wire_w_lg_w_lg_end_operation422w423w(0) <= wire_w_lg_end_operation422w(0) AND do_read_stat;
	wire_w_lg_w_lg_rden_wire315w316w(0) <= wire_w_lg_rden_wire315w(0) AND not_busy;
	wire_w_lg_do_4baddr150w(0) <= do_4baddr AND wire_w_lg_do_read_stat46w(0);
	wire_w_lg_do_bulk_erase254w(0) <= do_bulk_erase AND wire_w_lg_do_read_stat46w(0);
	wire_w_lg_do_polling420w(0) <= do_polling AND end_one_cyc_pos;
	wire_w_lg_do_sec_erase318w(0) <= do_sec_erase AND wire_w_lg_do_wren47w(0);
	wire_w_lg_do_sec_prot600w(0) <= do_sec_prot AND wire_spstage_cntr_w_lg_w_q_range598w599w(0);
	wire_w_lg_do_sec_prot612w(0) <= do_sec_prot AND stage3_wire;
	wire_w_lg_do_sec_prot621w(0) <= do_sec_prot AND wire_spstage_cntr_w_q_range598w(0);
	wire_w_lg_do_write171w(0) <= do_write AND wire_w_lg_do_read_stat46w(0);
	wire_w_lg_do_write63w(0) <= do_write AND wire_w_lg_w_pagewr_buf_not_empty_range61w62w(0);
	wire_w_lg_do_write56w(0) <= do_write AND shift_pgwr_data;
	wire_w_lg_end_operation409w(0) <= end_operation AND do_read_stat;
	wire_w_lg_load_opcode152w(0) <= load_opcode AND wire_w_lg_w_lg_do_4baddr150w151w(0);
	wire_w_lg_load_opcode173w(0) <= load_opcode AND wire_w_lg_w_lg_do_write171w172w(0);
	wire_w_lg_load_opcode158w(0) <= load_opcode AND do_bulk_erase;
	wire_w_lg_load_opcode176w(0) <= load_opcode AND do_fast_read;
	wire_w_lg_load_opcode179w(0) <= load_opcode AND do_read;
	wire_w_lg_load_opcode187w(0) <= load_opcode AND do_read_rdid;
	wire_w_lg_load_opcode190w(0) <= load_opcode AND do_read_sid;
	wire_w_lg_load_opcode168w(0) <= load_opcode AND do_read_stat;
	wire_w_lg_load_opcode163w(0) <= load_opcode AND do_sec_erase;
	wire_w_lg_load_opcode182w(0) <= load_opcode AND do_sec_prot;
	wire_w_lg_load_opcode155w(0) <= load_opcode AND do_wren;
	wire_w_lg_not_busy309w(0) <= not_busy AND wire_w_addr_range308w(0);
	loop12 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_not_busy304w(i) <= not_busy AND wire_w_addr_range303w(i);
	END GENERATE loop12;
	wire_w_lg_not_busy610w(0) <= not_busy AND wire_w_datain_range609w(0);
	loop13 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_not_busy605w(i) <= not_busy AND wire_w_datain_range604w(i);
	END GENERATE loop13;
	wire_w_lg_reach_max_cnt484w(0) <= reach_max_cnt AND shift_bytes_wire;
	wire_w_lg_read_bufdly447w(0) <= read_bufdly AND wire_scfifo4_w_q_range446w(0);
	loop14 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_read_bufdly442w(i) <= read_bufdly AND wire_scfifo4_w_q_range441w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_shift_opcode148w(i) <= shift_opcode AND wire_asmi_opcode_reg_w_q_range147w(i);
	END GENERATE loop15;
	wire_w_lg_stage3_wire314w(0) <= stage3_wire AND wire_w_lg_w_lg_w_lg_w_lg_do_write65w311w312w313w(0);
	wire_w_lg_stage3_wire341w(0) <= stage3_wire AND wire_w_lg_do_read_stat340w(0);
	loop16 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_stage3_wire302w(i) <= stage3_wire AND wire_addr_reg_w_q_range301w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_stage3_wire603w(i) <= stage3_wire AND wire_wrstat_dreg_w_q_range602w(i);
	END GENERATE loop17;
	wire_w_lg_stage4_wire343w(0) <= stage4_wire AND wire_w_lg_w_lg_do_read330w342w(0);
	wire_w_lg_start_poll259w(0) <= start_poll AND do_read_stat;
	wire_w_lg_wren_wire615w(0) <= wren_wire AND not_busy;
	wire_w_lg_w_lg_do_write56w272w(0) <= NOT wire_w_lg_do_write56w(0);
	wire_w_lg_bp0_wire516w(0) <= NOT bp0_wire;
	wire_w_lg_bp1_wire511w(0) <= NOT bp1_wire;
	wire_w_lg_bp2_wire522w(0) <= NOT bp2_wire;
	wire_w_lg_buf_empty553w(0) <= NOT buf_empty;
	wire_w_lg_busy_wire2w(0) <= NOT busy_wire;
	wire_w_lg_clkin_wire42w(0) <= NOT clkin_wire;
	wire_w_lg_do_4baddr404w(0) <= NOT do_4baddr;
	wire_w_lg_do_bulk_erase406w(0) <= NOT do_bulk_erase;
	wire_w_lg_do_fast_read273w(0) <= NOT do_fast_read;
	wire_w_lg_do_memadd327w(0) <= NOT do_memadd;
	wire_w_lg_do_polling268w(0) <= NOT do_polling;
	wire_w_lg_do_read274w(0) <= NOT do_read;
	wire_w_lg_do_read_rdid45w(0) <= NOT do_read_rdid;
	wire_w_lg_do_read_stat46w(0) <= NOT do_read_stat;
	wire_w_lg_do_sec_erase407w(0) <= NOT do_sec_erase;
	wire_w_lg_do_sec_prot405w(0) <= NOT do_sec_prot;
	wire_w_lg_do_wren47w(0) <= NOT do_wren;
	wire_w_lg_do_write408w(0) <= NOT do_write;
	wire_w_lg_end_add_cycle75w(0) <= NOT end_add_cycle;
	wire_w_lg_end_fast_read69w(0) <= NOT end_fast_read;
	wire_w_lg_end_ophdly43w(0) <= NOT end_ophdly;
	wire_w_lg_end_pgwr_data55w(0) <= NOT end_pgwr_data;
	wire_w_lg_end_read72w(0) <= NOT end_read;
	wire_w_lg_rden_wire389w(0) <= NOT rden_wire;
	wire_w_lg_reach_max_cnt449w(0) <= NOT reach_max_cnt;
	wire_w_lg_read_bufdly439w(0) <= NOT read_bufdly;
	wire_w_lg_read_rdid_wire11w(0) <= NOT read_rdid_wire;
	wire_w_lg_read_sid_wire10w(0) <= NOT read_sid_wire;
	wire_w_lg_read_status_wire26w(0) <= NOT read_status_wire;
	wire_w_lg_sec_erase_wire29w(0) <= NOT sec_erase_wire;
	wire_w_lg_sec_protect_wire14w(0) <= NOT sec_protect_wire;
	wire_w_lg_st_busy_wire102w(0) <= NOT st_busy_wire;
	wire_w_lg_write_prot_true487w(0) <= NOT write_prot_true;
	wire_w_lg_write_wire21w(0) <= NOT write_wire;
	wire_w_lg_w_pagewr_buf_not_empty_range61w62w(0) <= NOT wire_w_pagewr_buf_not_empty_range61w(0);
	wire_w_lg_w_lg_w586w587w588w(0) <= wire_w_lg_w586w587w(0) OR write_prot_true;
	wire_w_lg_w_lg_w_lg_load_opcode190w226w227w(0) <= wire_w_lg_w_lg_load_opcode190w226w(0) OR wire_w_lg_w_lg_load_opcode187w224w(0);
	loop18 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode190w191w192w(i) <= wire_w_lg_w_lg_load_opcode190w191w(i) OR wire_w_lg_w_lg_load_opcode187w188w(i);
	END GENERATE loop18;
	wire_w_lg_w_lg_w_lg_w_lg_do_write65w66w488w489w(0) <= wire_w_lg_w_lg_w_lg_do_write65w66w488w(0) OR do_4baddr;
	wire_w_lg_w_lg_w_lg_do_write65w311w312w(0) <= wire_w_lg_w_lg_do_write65w311w(0) OR do_read;
	wire_w_lg_w_lg_w_lg_rden_wire315w316w317w(0) <= wire_w_lg_w_lg_rden_wire315w316w(0) OR wire_w_lg_stage3_wire314w(0);
	loop19 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_not_busy304w305w(i) <= wire_w_lg_not_busy304w(i) OR wire_w_lg_stage3_wire302w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_not_busy605w606w(i) <= wire_w_lg_not_busy605w(i) OR wire_w_lg_stage3_wire603w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_read_bufdly442w443w(i) <= wire_w_lg_read_bufdly442w(i) OR wire_w_lg_w_lg_read_bufdly439w440w(i);
	END GENERATE loop21;
	wire_w_lg_w_lg_stage4_wire343w344w(0) <= wire_w_lg_stage4_wire343w(0) OR wire_w_lg_stage3_wire341w(0);
	wire_w_lg_w_lg_wren_wire615w616w(0) <= wire_w_lg_wren_wire615w(0) OR wire_w_lg_w_lg_w_lg_do_sec_prot612w613w614w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode190w226w227w228w(0) <= wire_w_lg_w_lg_w_lg_load_opcode190w226w227w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode182w183w184w222w(0);
	loop22 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode190w191w192w193w(i) <= wire_w_lg_w_lg_w_lg_load_opcode190w191w192w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode182w183w184w185w(i);
	END GENERATE loop22;
	wire_w_lg_w_lg_w_lg_w_lg_do_write65w311w312w313w(0) <= wire_w_lg_w_lg_w_lg_do_write65w311w312w(0) OR do_fast_read;
	wire_w229w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode190w226w227w228w(0) OR wire_w_lg_w_lg_load_opcode179w220w(0);
	loop23 : FOR i IN 0 TO 6 GENERATE 
		wire_w194w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode190w191w192w193w(i) OR wire_w_lg_w_lg_load_opcode179w180w(i);
	END GENERATE loop23;
	wire_w_lg_w229w230w(0) <= wire_w229w(0) OR wire_w_lg_w_lg_load_opcode176w218w(0);
	loop24 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w194w195w(i) <= wire_w194w(i) OR wire_w_lg_w_lg_load_opcode176w177w(i);
	END GENERATE loop24;
	wire_w_lg_w_lg_w229w230w231w(0) <= wire_w_lg_w229w230w(0) OR wire_w_lg_w_lg_load_opcode173w216w(0);
	loop25 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w194w195w196w(i) <= wire_w_lg_w194w195w(i) OR wire_w_lg_w_lg_load_opcode173w174w(i);
	END GENERATE loop25;
	wire_w_lg_w_lg_w_lg_w229w230w231w232w(0) <= wire_w_lg_w_lg_w229w230w231w(0) OR wire_w_lg_w_lg_load_opcode168w214w(0);
	loop26 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w194w195w196w197w(i) <= wire_w_lg_w_lg_w194w195w196w(i) OR wire_w_lg_w_lg_load_opcode168w169w(i);
	END GENERATE loop26;
	wire_w_lg_w_lg_w_lg_w_lg_w229w230w231w232w233w(0) <= wire_w_lg_w_lg_w_lg_w229w230w231w232w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode163w164w165w212w(0);
	loop27 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w194w195w196w197w198w(i) <= wire_w_lg_w_lg_w_lg_w194w195w196w197w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode163w164w165w166w(i);
	END GENERATE loop27;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w229w230w231w232w233w234w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w229w230w231w232w233w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode158w159w160w210w(0);
	loop28 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w_lg_w194w195w196w197w198w199w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w194w195w196w197w198w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode158w159w160w161w(i);
	END GENERATE loop28;
	wire_w235w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w229w230w231w232w233w234w(0) OR wire_w_lg_w_lg_load_opcode155w208w(0);
	loop29 : FOR i IN 0 TO 6 GENERATE 
		wire_w200w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w194w195w196w197w198w199w(i) OR wire_w_lg_w_lg_load_opcode155w156w(i);
	END GENERATE loop29;
	wire_w_lg_w235w236w(0) <= wire_w235w(0) OR wire_w_lg_w_lg_load_opcode152w206w(0);
	loop30 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w200w201w(i) <= wire_w200w(i) OR wire_w_lg_w_lg_load_opcode152w153w(i);
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w200w201w202w(i) <= wire_w_lg_w200w201w(i) OR wire_w_lg_shift_opcode148w(i);
	END GENERATE loop31;
	wire_w134w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read_sid130w131w132w133w(0) OR do_read_rdid;
	wire_w_lg_w_lg_w_lg_w_lg_do_read_sid130w131w132w133w(0) <= wire_w_lg_w_lg_w_lg_do_read_sid130w131w132w(0) OR do_sec_erase;
	wire_w_lg_w_lg_w_lg_do_read330w331w332w(0) <= wire_w_lg_w_lg_do_read330w331w(0) OR do_sec_erase;
	wire_w_lg_w_lg_w_lg_do_read_sid130w131w132w(0) <= wire_w_lg_w_lg_do_read_sid130w131w(0) OR do_write;
	wire_w_lg_w_lg_w_lg_do_write65w66w499w(0) <= wire_w_lg_w_lg_do_write65w66w(0) OR do_4baddr;
	wire_w_lg_w_lg_do_read330w342w(0) <= wire_w_lg_do_read330w(0) OR do_read_sid;
	wire_w_lg_w_lg_do_read330w331w(0) <= wire_w_lg_do_read330w(0) OR do_write;
	wire_w_lg_w_lg_do_read_sid130w131w(0) <= wire_w_lg_do_read_sid130w(0) OR do_fast_read;
	wire_w_lg_w_lg_do_sec_erase501w502w(0) <= wire_w_lg_do_sec_erase501w(0) OR do_bulk_erase;
	wire_w_lg_w_lg_do_write65w66w(0) <= wire_w_lg_do_write65w(0) OR do_bulk_erase;
	wire_w_lg_data0out_wire346w(0) <= data0out_wire OR wire_w_dataout_wire_range345w(0);
	wire_w_lg_do_4baddr255w(0) <= do_4baddr OR wire_w_lg_do_bulk_erase254w(0);
	wire_w_lg_do_read330w(0) <= do_read OR do_fast_read;
	wire_w_lg_do_read_sid130w(0) <= do_read_sid OR do_read;
	wire_w_lg_do_read_stat340w(0) <= do_read_stat OR do_read_rdid;
	wire_w_lg_do_sec_erase501w(0) <= do_sec_erase OR do_write;
	wire_w_lg_do_wren256w(0) <= do_wren OR wire_w_lg_do_4baddr255w(0);
	wire_w_lg_do_write65w(0) <= do_write OR do_sec_erase;
	wire_w_lg_end_operation422w(0) <= end_operation OR wire_w_lg_w_lg_do_polling420w421w(0);
	wire_w_lg_load_opcode238w(0) <= load_opcode OR shift_opcode;
	wire_w_lg_rden_wire315w(0) <= rden_wire OR wren_wire;
	wire_w_lg_read_bufdly437w(0) <= read_bufdly OR shift_pgwr_data;
	wire_w_lg_w_pagewr_buf_not_empty_range453w456w(0) <= wire_w_pagewr_buf_not_empty_range453w(0) OR wire_pgwr_data_cntr_w_q_range455w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range457w459w(0) <= wire_w_pagewr_buf_not_empty_range457w(0) OR wire_pgwr_data_cntr_w_q_range458w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range460w462w(0) <= wire_w_pagewr_buf_not_empty_range460w(0) OR wire_pgwr_data_cntr_w_q_range461w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range463w465w(0) <= wire_w_pagewr_buf_not_empty_range463w(0) OR wire_pgwr_data_cntr_w_q_range464w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range466w468w(0) <= wire_w_pagewr_buf_not_empty_range466w(0) OR wire_pgwr_data_cntr_w_q_range467w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range469w471w(0) <= wire_w_pagewr_buf_not_empty_range469w(0) OR wire_pgwr_data_cntr_w_q_range470w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range472w474w(0) <= wire_w_pagewr_buf_not_empty_range472w(0) OR wire_pgwr_data_cntr_w_q_range473w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range475w477w(0) <= wire_w_pagewr_buf_not_empty_range475w(0) OR wire_pgwr_data_cntr_w_q_range476w(0);
	b4addr_opcode <= (OTHERS => '0');
	be_write_prot <= (do_bulk_erase AND (((bp3_wire OR bp2_wire) OR bp1_wire) OR bp0_wire));
	berase_opcode <= "11000111";
	bp0_wire <= statreg_int(2);
	bp1_wire <= statreg_int(3);
	bp2_wire <= statreg_int(4);
	bp3_wire <= statreg_int(6);
	buf_empty <= buf_empty_reg;
	bulk_erase_wire <= bulk_erase_reg;
	busy <= (busy_wire OR busy_delay_reg);
	busy_wire <= (((((((((do_read_rdid OR do_read_sid) OR do_read) OR do_fast_read) OR do_write) OR do_sec_prot) OR do_read_stat) OR do_sec_erase) OR do_bulk_erase) OR do_4baddr);
	clkin_wire <= clkin;
	clr_rdid_wire <= clr_rdid_reg2;
	clr_read_wire <= clr_read_reg2;
	clr_rstat_wire <= clr_rstat_reg2;
	clr_secprot_wire <= clr_secprot_reg2;
	clr_write_wire <= clr_write_reg2;
	cnt_bfend_wire_in <= (wire_gen_cntr_w_lg_w_q_range99w100w(0) AND wire_gen_cntr_q(0));
	data0out_wire <= wire_cycloneii_asmiblock3_data0out;
	data_valid <= data_valid_wire;
	data_valid_wire <= dvalid_reg2;
	dataout <= ( read_data_reg(7 DOWNTO 0));
	dataout_wire <= ( "0000");
	do_4baddr <= '0';
	do_bulk_erase <= (((((((wire_w_lg_read_rdid_wire11w(0) AND wire_w_lg_read_sid_wire10w(0)) AND wire_w_lg_sec_protect_wire14w(0)) AND (NOT (read_wire OR fast_read_wire))) AND wire_w_lg_write_wire21w(0)) AND wire_w_lg_read_status_wire26w(0)) AND wire_w_lg_sec_erase_wire29w(0)) AND bulk_erase_wire);
	do_fast_read <= (((wire_w_lg_read_rdid_wire11w(0) AND wire_w_lg_read_sid_wire10w(0)) AND wire_w_lg_sec_protect_wire14w(0)) AND fast_read_wire);
	do_memadd <= do_wrmemadd_reg;
	do_polling <= (do_write_polling OR do_sprot_polling);
	do_read <= '0';
	do_read_rdid <= read_rdid_wire;
	do_read_sid <= '0';
	do_read_stat <= (((((((wire_w_lg_read_rdid_wire11w(0) AND wire_w_lg_read_sid_wire10w(0)) AND wire_w_lg_sec_protect_wire14w(0)) AND (NOT (read_wire OR fast_read_wire))) AND wire_w_lg_write_wire21w(0)) AND read_status_wire) OR do_write_rstat) OR do_sprot_rstat);
	do_sec_erase <= ((((((wire_w_lg_read_rdid_wire11w(0) AND wire_w_lg_read_sid_wire10w(0)) AND wire_w_lg_sec_protect_wire14w(0)) AND (NOT (read_wire OR fast_read_wire))) AND wire_w_lg_write_wire21w(0)) AND wire_w_lg_read_status_wire26w(0)) AND sec_erase_wire);
	do_sec_prot <= ((wire_w_lg_read_rdid_wire11w(0) AND wire_w_lg_read_sid_wire10w(0)) AND sec_protect_wire);
	do_secprot_wren <= (wire_w_lg_do_sec_prot600w(0) AND (NOT wire_spstage_cntr_q(0)));
	do_sprot_polling <= (wire_w_lg_do_sec_prot621w(0) AND wire_spstage_cntr_q(0));
	do_sprot_rstat <= sprot_rstat_reg;
	do_wren <= (do_write_wren OR do_secprot_wren);
	do_write <= ((((wire_w_lg_read_rdid_wire11w(0) AND wire_w_lg_read_sid_wire10w(0)) AND wire_w_lg_sec_protect_wire14w(0)) AND (NOT (read_wire OR fast_read_wire))) AND write_wire);
	do_write_polling <= ((wire_w_lg_w_lg_do_write65w66w(0) AND wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_w_lg_w_q_range492w493w(0));
	do_write_rstat <= write_rstat_reg;
	do_write_wren <= ((NOT wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_q(0));
	dummy_read_buf <= maxcnt_shift_reg2;
	end1_cyc_dlyncs_in_wire <= (((((((((wire_stage_cntr_w_lg_w_lg_w_q_range88w93w107w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND (NOT wire_gen_cntr_q(0))) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w93w107w108w109w(0)) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read)) OR wire_w_lg_w_lg_w_lg_do_write65w66w67w(0)) OR wire_w_lg_do_write63w(0)) OR ((do_read_stat AND start_poll) AND wire_w_lg_st_busy_wire102w(0)));
	end1_cyc_gen_cntr_wire <= (wire_gen_cntr_w_lg_w_q_range99w100w(0) AND (NOT wire_gen_cntr_q(0)));
	end1_cyc_normal_in_wire <= (((((((((wire_stage_cntr_w_lg_w_lg_w_q_range88w93w107w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND wire_gen_cntr_q(0)) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w93w107w108w109w(0)) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read)) OR wire_w_lg_w_lg_w_lg_do_write65w66w67w(0)) OR wire_w_lg_do_write63w(0)) OR ((do_read_stat AND start_poll) AND wire_w_lg_st_busy_wire102w(0)));
	end1_cyc_reg_in_wire <= wire_mux211_dataout;
	end_add_cycle <= wire_mux212_dataout;
	end_add_cycle_mux_datab_wire <= (wire_addbyte_cntr_q(2) AND wire_addbyte_cntr_q(1));
	end_fast_read <= end_read_reg;
	end_one_cyc_pos <= end1_cyc_reg2;
	end_one_cycle <= end1_cyc_reg;
	end_operation <= end_op_reg;
	end_opfdly <= end_opfdly_reg;
	end_ophdly <= end_op_hdlyreg;
	end_pgwr_data <= end_pgwrop_reg;
	end_read <= end_read_reg;
	end_read_byte <= end_rbyte_reg;
	end_wrstage <= end_operation;
	fast_read_opcode <= "00001011";
	fast_read_wire <= fast_read_reg;
	ill_erase_wire <= ill_erase_reg;
	ill_write_wire <= ill_write_reg;
	illegal_erase <= ill_erase_wire;
	illegal_erase_b4out_wire <= ((do_sec_erase OR do_bulk_erase) AND write_prot_true);
	illegal_write <= ill_write_wire;
	illegal_write_b4out_wire <= ((do_write AND write_prot_true) OR wire_w_lg_do_write63w(0));
	in_operation <= busy_wire;
	load_opcode <= ((((wire_stage_cntr_w_lg_w_q_range89w90w(0) AND wire_stage_cntr_w_lg_w_q_range88w93w(0)) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_w_lg_w_q_range97w98w(0)) AND wire_gen_cntr_q(0));
	memadd_sdoin <= add_msb_reg;
	not_busy <= busy_det_reg;
	oe_wire <= '0';
	page_size_wire <= "100000000";
	pagewr_buf_not_empty <= ( wire_w_lg_w_pagewr_buf_not_empty_range475w477w & wire_w_lg_w_pagewr_buf_not_empty_range472w474w & wire_w_lg_w_pagewr_buf_not_empty_range469w471w & wire_w_lg_w_pagewr_buf_not_empty_range466w468w & wire_w_lg_w_pagewr_buf_not_empty_range463w465w & wire_w_lg_w_pagewr_buf_not_empty_range460w462w & wire_w_lg_w_pagewr_buf_not_empty_range457w459w & wire_w_lg_w_pagewr_buf_not_empty_range453w456w & wire_pgwr_data_cntr_q(0));
	rden_wire <= rden;
	rdid_load <= (end_operation AND do_read_rdid);
	rdid_opcode <= "10011111";
	rdid_out <= ( rdid_out_reg(7 DOWNTO 0));
	reach_max_cnt <= max_cnt_reg;
	read_buf <= (((((end_one_cycle AND do_write) AND wire_w_lg_do_read_stat46w(0)) AND wire_w_lg_do_wren47w(0)) AND (wire_stage_cntr_w_lg_w_q_range89w94w(0) OR wire_addbyte_cntr_w_lg_w_q_range137w142w(0))) AND wire_w_lg_buf_empty553w(0));
	read_bufdly <= read_bufdly_reg;
	read_data_reg_in_wire <= ( read_dout_reg(7 DOWNTO 0));
	read_opcode <= (OTHERS => '0');
	read_rdid_wire <= read_rdid_reg;
	read_sid_wire <= '0';
	read_status_wire <= read_status_reg;
	read_wire <= '0';
	rsid_opcode <= (OTHERS => '0');
	rsid_sdoin <= '0';
	rstat_opcode <= "00000101";
	scein_wire <= wire_ncs_reg_w_lg_q291w(0);
	sdoin_wire <= to_sdoin_wire;
	sec_erase_wire <= sec_erase_reg;
	sec_protect_wire <= sec_prot_reg;
	secprot_opcode <= "00000001";
	secprot_sdoin <= (stage3_wire AND streg_datain_reg);
	serase_opcode <= "11011000";
	shift_bytes_wire <= shift_bytes;
	shift_opcode <= shift_op_reg;
	shift_opdata <= stage2_wire;
	shift_pgwr_data <= shftpgwr_data_reg;
	st_busy_wire <= statreg_int(0);
	stage2_wire <= stage2_reg;
	stage3_wire <= stage3_reg;
	stage4_wire <= stage4_reg;
	start_poll <= (start_wrpoll OR start_sppoll);
	start_sppoll <= start_sppoll_reg2;
	start_wrpoll <= start_wrpoll_reg2;
	status_out <= ( statreg_out(7 DOWNTO 0));
	to_sdoin_wire <= (((((shift_opdata AND asmi_opcode_reg(7)) OR rsid_sdoin) OR memadd_sdoin) OR write_sdoin) OR secprot_sdoin);
	wren_opcode <= "00000110";
	wren_wire <= wren;
	write_opcode <= "00000010";
	write_prot_true <= write_prot_reg;
	write_sdoin <= ((((do_write AND stage4_wire) AND wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_q(0)) AND pgwrbuf_dataout(7));
	write_wire <= write_reg;
	wire_w_addr_range308w(0) <= addr(0);
	wire_w_addr_range303w <= addr(23 DOWNTO 1);
	wire_w_b4addr_opcode_range205w(0) <= b4addr_opcode(0);
	wire_w_b4addr_opcode_range149w <= b4addr_opcode(7 DOWNTO 1);
	wire_w_berase_opcode_range209w(0) <= berase_opcode(0);
	wire_w_berase_opcode_range157w <= berase_opcode(7 DOWNTO 1);
	wire_w_datain_range609w(0) <= datain(0);
	wire_w_datain_range604w <= datain(7 DOWNTO 1);
	wire_w_dataout_wire_range345w(0) <= dataout_wire(1);
	wire_w_fast_read_opcode_range217w(0) <= fast_read_opcode(0);
	wire_w_fast_read_opcode_range175w <= fast_read_opcode(7 DOWNTO 1);
	wire_w_pagewr_buf_not_empty_range453w(0) <= pagewr_buf_not_empty(0);
	wire_w_pagewr_buf_not_empty_range457w(0) <= pagewr_buf_not_empty(1);
	wire_w_pagewr_buf_not_empty_range460w(0) <= pagewr_buf_not_empty(2);
	wire_w_pagewr_buf_not_empty_range463w(0) <= pagewr_buf_not_empty(3);
	wire_w_pagewr_buf_not_empty_range466w(0) <= pagewr_buf_not_empty(4);
	wire_w_pagewr_buf_not_empty_range469w(0) <= pagewr_buf_not_empty(5);
	wire_w_pagewr_buf_not_empty_range472w(0) <= pagewr_buf_not_empty(6);
	wire_w_pagewr_buf_not_empty_range475w(0) <= pagewr_buf_not_empty(7);
	wire_w_pagewr_buf_not_empty_range61w(0) <= pagewr_buf_not_empty(8);
	wire_w_rdid_opcode_range223w(0) <= rdid_opcode(0);
	wire_w_rdid_opcode_range186w <= rdid_opcode(7 DOWNTO 1);
	wire_w_read_opcode_range219w(0) <= read_opcode(0);
	wire_w_read_opcode_range178w <= read_opcode(7 DOWNTO 1);
	wire_w_rsid_opcode_range225w(0) <= rsid_opcode(0);
	wire_w_rsid_opcode_range189w <= rsid_opcode(7 DOWNTO 1);
	wire_w_rstat_opcode_range213w(0) <= rstat_opcode(0);
	wire_w_rstat_opcode_range167w <= rstat_opcode(7 DOWNTO 1);
	wire_w_secprot_opcode_range221w(0) <= secprot_opcode(0);
	wire_w_secprot_opcode_range181w <= secprot_opcode(7 DOWNTO 1);
	wire_w_serase_opcode_range211w(0) <= serase_opcode(0);
	wire_w_serase_opcode_range162w <= serase_opcode(7 DOWNTO 1);
	wire_w_wren_opcode_range207w(0) <= wren_opcode(0);
	wire_w_wren_opcode_range154w <= wren_opcode(7 DOWNTO 1);
	wire_w_write_opcode_range215w(0) <= write_opcode(0);
	wire_w_write_opcode_range170w <= write_opcode(7 DOWNTO 1);
	wire_addbyte_cntr_w_lg_w_q_range137w142w(0) <= wire_addbyte_cntr_w_q_range137w(0) AND wire_addbyte_cntr_w_lg_w_q_range140w141w(0);
	wire_addbyte_cntr_w_lg_w_q_range140w141w(0) <= NOT wire_addbyte_cntr_w_q_range140w(0);
	wire_addbyte_cntr_clk_en <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w135w136w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w135w136w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range89w92w135w(0) AND wire_w134w(0);
	wire_addbyte_cntr_clock <= wire_w_lg_clkin_wire42w(0);
	wire_addbyte_cntr_w_q_range140w(0) <= wire_addbyte_cntr_q(0);
	wire_addbyte_cntr_w_q_range137w(0) <= wire_addbyte_cntr_q(1);
	addbyte_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => end_operation,
		clk_en => wire_addbyte_cntr_clk_en,
		clock => wire_addbyte_cntr_clock,
		q => wire_addbyte_cntr_q
	  );
	wire_gen_cntr_w_lg_w_q_range99w100w(0) <= wire_gen_cntr_w_q_range99w(0) AND wire_gen_cntr_w_lg_w_q_range97w98w(0);
	wire_gen_cntr_w_lg_w_q_range97w98w(0) <= NOT wire_gen_cntr_w_q_range97w(0);
	wire_gen_cntr_clk_en <= wire_w_lg_in_operation44w(0);
	wire_w_lg_in_operation44w(0) <= in_operation AND wire_w_lg_end_ophdly43w(0);
	wire_gen_cntr_w_q_range97w(0) <= wire_gen_cntr_q(1);
	wire_gen_cntr_w_q_range99w(0) <= wire_gen_cntr_q(2);
	gen_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => end_one_cycle,
		clk_en => wire_gen_cntr_clk_en,
		clock => clkin_wire,
		q => wire_gen_cntr_q
	  );
	wire_spstage_cntr_w_lg_w_q_range598w599w(0) <= NOT wire_spstage_cntr_w_q_range598w(0);
	wire_spstage_cntr_clk_en <= wire_w_lg_do_sec_prot595w(0);
	wire_w_lg_do_sec_prot595w(0) <= do_sec_prot AND end_operation;
	wire_spstage_cntr_clock <= wire_w_lg_clkin_wire42w(0);
	wire_spstage_cntr_w_q_range596w(0) <= wire_spstage_cntr_q(0);
	wire_spstage_cntr_w_q_range598w(0) <= wire_spstage_cntr_q(1);
	spstage_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 2
	  )
	  PORT MAP ( 
		aclr => clr_secprot_wire,
		clk_en => wire_spstage_cntr_clk_en,
		clock => wire_spstage_cntr_clock,
		q => wire_spstage_cntr_q
	  );
	wire_stage_cntr_w_lg_w247w248w(0) <= wire_stage_cntr_w247w(0) AND end_one_cycle;
	wire_stage_cntr_w247w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w92w244w245w246w(0) AND end_add_cycle;
	wire_stage_cntr_w252w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w92w249w250w251w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w92w244w245w246w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w244w245w(0) AND wire_w_lg_do_read_stat46w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w92w249w250w251w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w249w250w(0) AND wire_w_lg_do_read_stat46w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w90w91w257w258w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w90w91w257w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w94w322w323w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range89w94w322w(0) AND end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w269w270w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range89w92w269w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w244w245w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range89w92w244w(0) AND wire_w_lg_do_wren47w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w249w250w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range89w92w249w(0) AND wire_w_lg_do_wren47w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w90w91w257w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range89w90w91w(0) AND wire_w_lg_do_wren256w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range89w94w322w(0) <= wire_stage_cntr_w_lg_w_q_range89w94w(0) AND end_add_cycle;
	wire_stage_cntr_w_lg_w_lg_w_q_range89w92w269w(0) <= wire_stage_cntr_w_lg_w_q_range89w92w(0) AND do_read_stat;
	wire_stage_cntr_w_lg_w_lg_w_q_range89w92w244w(0) <= wire_stage_cntr_w_lg_w_q_range89w92w(0) AND do_sec_erase;
	wire_stage_cntr_w_lg_w_lg_w_q_range89w92w249w(0) <= wire_stage_cntr_w_lg_w_q_range89w92w(0) AND do_sec_prot;
	wire_stage_cntr_w_lg_w_lg_w_q_range89w92w135w(0) <= wire_stage_cntr_w_lg_w_q_range89w92w(0) AND end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w93w107w108w109w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w93w107w108w(0) AND end1_cyc_gen_cntr_wire;
	wire_stage_cntr_w_lg_w_lg_w_q_range88w93w107w(0) <= wire_stage_cntr_w_lg_w_q_range88w93w(0) AND wire_stage_cntr_w_lg_w_q_range89w90w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range89w90w91w(0) <= wire_stage_cntr_w_lg_w_q_range89w90w(0) AND wire_stage_cntr_w_q_range88w(0);
	wire_stage_cntr_w_lg_w_q_range89w94w(0) <= wire_stage_cntr_w_q_range89w(0) AND wire_stage_cntr_w_lg_w_q_range88w93w(0);
	wire_stage_cntr_w_lg_w_q_range89w92w(0) <= wire_stage_cntr_w_q_range89w(0) AND wire_stage_cntr_w_q_range88w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w93w107w108w(0) <= NOT wire_stage_cntr_w_lg_w_lg_w_q_range88w93w107w(0);
	wire_stage_cntr_w_lg_w_q_range88w93w(0) <= NOT wire_stage_cntr_w_q_range88w(0);
	wire_stage_cntr_w_lg_w_q_range89w90w(0) <= NOT wire_stage_cntr_w_q_range89w(0);
	wire_stage_cntr_clk_en <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w82w83w84w85w86w87w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w82w83w84w85w86w87w(0) <= (((((((((in_operation AND end_one_cycle) AND (NOT (stage3_wire AND wire_w_lg_end_add_cycle75w(0)))) AND (NOT (stage4_wire AND wire_w_lg_end_read72w(0)))) AND (NOT (stage4_wire AND wire_w_lg_end_fast_read69w(0)))) AND (NOT wire_w_lg_w_lg_w_lg_do_write65w66w67w(0))) AND (NOT wire_w_lg_do_write63w(0))) AND (NOT (stage3_wire AND st_busy_wire))) AND (NOT (wire_w_lg_do_write56w(0) AND wire_w_lg_end_pgwr_data55w(0)))) AND (NOT (stage2_wire AND do_wren))) AND (NOT ((((stage3_wire AND do_sec_erase) AND wire_w_lg_do_wren47w(0)) AND wire_w_lg_do_read_stat46w(0)) AND wire_w_lg_do_read_rdid45w(0)));
	wire_stage_cntr_w_q_range88w(0) <= wire_stage_cntr_q(0);
	wire_stage_cntr_w_q_range89w(0) <= wire_stage_cntr_q(1);
	stage_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 2
	  )
	  PORT MAP ( 
		aclr => end_ophdly,
		clk_en => wire_stage_cntr_clk_en,
		clock => clkin_wire,
		q => wire_stage_cntr_q
	  );
	wire_wrstage_cntr_w_lg_w_q_range494w495w(0) <= wire_wrstage_cntr_w_q_range494w(0) AND wire_wrstage_cntr_w_lg_w_q_range492w493w(0);
	wire_wrstage_cntr_w_lg_w_q_range492w493w(0) <= NOT wire_wrstage_cntr_w_q_range492w(0);
	wire_wrstage_cntr_clk_en <= wire_w_lg_w490w491w(0);
	wire_w_lg_w490w491w(0) <= wire_w490w(0) AND wire_w_lg_st_busy_wire102w(0);
	wire_wrstage_cntr_clock <= wire_w_lg_clkin_wire42w(0);
	wire_wrstage_cntr_w_q_range492w(0) <= wire_wrstage_cntr_q(0);
	wire_wrstage_cntr_w_q_range494w(0) <= wire_wrstage_cntr_q(1);
	wrstage_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 2
	  )
	  PORT MAP ( 
		aclr => clr_write_wire,
		clk_en => wire_wrstage_cntr_clk_en,
		clock => wire_wrstage_cntr_clock,
		q => wire_wrstage_cntr_q
	  );
	cycloneii_asmiblock3 :  cycloneii_asmiblock
	  PORT MAP ( 
		data0out => wire_cycloneii_asmiblock3_data0out,
		dclkin => clkin_wire,
		oe => oe_wire,
		scein => scein_wire,
		sdoin => sdoin_wire
	  );
	PROCESS (clkin_wire, clr_addmsb_reg)
	BEGIN
		IF (clr_addmsb_reg = '1') THEN add_msb_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_add_msb_reg_ena = '1') THEN add_msb_reg <= addr_reg(23);
			END IF;
		END IF;
	END PROCESS;
	wire_add_msb_reg_ena <= (((wire_w_lg_w_lg_w_lg_do_read330w331w332w(0) AND (NOT (wire_w_lg_do_write65w(0) AND wire_w_lg_do_memadd327w(0)))) AND wire_stage_cntr_q(1)) AND wire_stage_cntr_q(0));
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(0) = '1') THEN addr_reg(0) <= wire_addr_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(1) = '1') THEN addr_reg(1) <= wire_addr_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(2) = '1') THEN addr_reg(2) <= wire_addr_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(3) = '1') THEN addr_reg(3) <= wire_addr_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(4) = '1') THEN addr_reg(4) <= wire_addr_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(5) = '1') THEN addr_reg(5) <= wire_addr_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(6) = '1') THEN addr_reg(6) <= wire_addr_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(7) = '1') THEN addr_reg(7) <= wire_addr_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(8) = '1') THEN addr_reg(8) <= wire_addr_reg_d(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(9) = '1') THEN addr_reg(9) <= wire_addr_reg_d(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(10) = '1') THEN addr_reg(10) <= wire_addr_reg_d(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(11) = '1') THEN addr_reg(11) <= wire_addr_reg_d(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(12) = '1') THEN addr_reg(12) <= wire_addr_reg_d(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(13) = '1') THEN addr_reg(13) <= wire_addr_reg_d(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(14) = '1') THEN addr_reg(14) <= wire_addr_reg_d(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(15) = '1') THEN addr_reg(15) <= wire_addr_reg_d(15);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(16) = '1') THEN addr_reg(16) <= wire_addr_reg_d(16);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(17) = '1') THEN addr_reg(17) <= wire_addr_reg_d(17);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(18) = '1') THEN addr_reg(18) <= wire_addr_reg_d(18);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(19) = '1') THEN addr_reg(19) <= wire_addr_reg_d(19);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(20) = '1') THEN addr_reg(20) <= wire_addr_reg_d(20);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(21) = '1') THEN addr_reg(21) <= wire_addr_reg_d(21);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(22) = '1') THEN addr_reg(22) <= wire_addr_reg_d(22);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(23) = '1') THEN addr_reg(23) <= wire_addr_reg_d(23);
			END IF;
		END IF;
	END PROCESS;
	wire_addr_reg_d <= ( wire_w_lg_w_lg_not_busy304w305w & wire_w_lg_not_busy309w);
	loop32 : FOR i IN 0 TO 23 GENERATE
		wire_addr_reg_ena(i) <= wire_w_lg_w_lg_w_lg_rden_wire315w316w317w(0);
	END GENERATE loop32;
	wire_addr_reg_w_lg_w_lg_w535w536w537w(0) <= wire_addr_reg_w_lg_w535w536w(0) AND bp0_wire;
	wire_addr_reg_w_lg_w535w536w(0) <= wire_addr_reg_w535w(0) AND wire_w_lg_bp1_wire511w(0);
	wire_addr_reg_w527w(0) <= wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range512w518w524w525w526w(0) AND bp0_wire;
	wire_addr_reg_w531w(0) <= wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range512w518w524w529w530w(0) AND bp1_wire;
	wire_addr_reg_w535w(0) <= wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range512w518w524w529w534w(0) AND wire_w_lg_bp2_wire522w(0);
	wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range512w518w524w525w526w(0) <= wire_addr_reg_w_lg_w_lg_w_lg_w_q_range512w518w524w525w(0) AND bp1_wire;
	wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range512w518w524w529w530w(0) <= wire_addr_reg_w_lg_w_lg_w_lg_w_q_range512w518w524w529w(0) AND wire_w_lg_bp2_wire522w(0);
	wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range512w518w524w529w534w(0) <= wire_addr_reg_w_lg_w_lg_w_lg_w_q_range512w518w524w529w(0) AND wire_addr_reg_w_q_range533w(0);
	wire_addr_reg_w_lg_w_lg_w_lg_w_q_range512w513w514w515w(0) <= wire_addr_reg_w_lg_w_lg_w_q_range512w513w514w(0) AND bp0_wire;
	wire_addr_reg_w_lg_w_lg_w_lg_w_q_range512w518w524w525w(0) <= wire_addr_reg_w_lg_w_lg_w_q_range512w518w524w(0) AND wire_w_lg_bp2_wire522w(0);
	wire_addr_reg_w_lg_w_lg_w_lg_w_q_range512w518w524w529w(0) <= wire_addr_reg_w_lg_w_lg_w_q_range512w518w524w(0) AND wire_addr_reg_w_q_range528w(0);
	wire_addr_reg_w_lg_w_lg_w_q_range512w513w514w(0) <= wire_addr_reg_w_lg_w_q_range512w513w(0) AND wire_w_lg_bp1_wire511w(0);
	wire_addr_reg_w_lg_w_lg_w_q_range512w518w519w(0) <= wire_addr_reg_w_lg_w_q_range512w518w(0) AND bp2_wire;
	wire_addr_reg_w_lg_w_lg_w_q_range512w518w524w(0) <= wire_addr_reg_w_lg_w_q_range512w518w(0) AND wire_addr_reg_w_q_range523w(0);
	wire_addr_reg_w_lg_w_q_range512w513w(0) <= wire_addr_reg_w_q_range512w(0) AND bp2_wire;
	wire_addr_reg_w_lg_w_q_range512w518w(0) <= wire_addr_reg_w_q_range512w(0) AND wire_addr_reg_w_q_range517w(0);
	wire_addr_reg_w_q_range533w(0) <= addr_reg(16);
	wire_addr_reg_w_q_range528w(0) <= addr_reg(17);
	wire_addr_reg_w_q_range523w(0) <= addr_reg(18);
	wire_addr_reg_w_q_range517w(0) <= addr_reg(19);
	wire_addr_reg_w_q_range512w(0) <= addr_reg(20);
	wire_addr_reg_w_q_range301w <= addr_reg(22 DOWNTO 0);
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(0) = '1') THEN asmi_opcode_reg(0) <= wire_asmi_opcode_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(1) = '1') THEN asmi_opcode_reg(1) <= wire_asmi_opcode_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(2) = '1') THEN asmi_opcode_reg(2) <= wire_asmi_opcode_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(3) = '1') THEN asmi_opcode_reg(3) <= wire_asmi_opcode_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(4) = '1') THEN asmi_opcode_reg(4) <= wire_asmi_opcode_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(5) = '1') THEN asmi_opcode_reg(5) <= wire_asmi_opcode_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(6) = '1') THEN asmi_opcode_reg(6) <= wire_asmi_opcode_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(7) = '1') THEN asmi_opcode_reg(7) <= wire_asmi_opcode_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_asmi_opcode_reg_d <= ( wire_w_lg_w_lg_w200w201w202w & wire_w_lg_w235w236w);
	loop33 : FOR i IN 0 TO 7 GENERATE
		wire_asmi_opcode_reg_ena(i) <= wire_w_lg_load_opcode238w(0);
	END GENERATE loop33;
	wire_asmi_opcode_reg_w_q_range147w <= asmi_opcode_reg(6 DOWNTO 0);
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN buf_empty_reg <= wire_cmpr6_aeb;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN bulk_erase_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_bulk_erase_reg_ena = '1') THEN bulk_erase_reg <= bulk_erase;
			END IF;
		END IF;
	END PROCESS;
	wire_bulk_erase_reg_ena <= (wire_w_lg_busy_wire2w(0) AND wren_wire);
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (power_up_reg = '1') THEN busy_delay_reg <= busy_wire;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN busy_det_reg <= wire_w_lg_busy_wire2w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_addmsb_reg <= ((wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w94w322w323w(0) OR wire_w_lg_w_lg_w_lg_do_read274w275w321w(0)) OR wire_w_lg_w_lg_w_lg_do_sec_erase318w319w320w(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN clr_endrbyte_reg <= ((((wire_w_lg_do_read330w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND wire_gen_cntr_q(0)) OR clr_read_wire);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_rdid_reg <= end_operation;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_rdid_reg2 <= clr_rdid_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_read_reg <= ((end_operation OR do_read_sid) OR do_sec_prot);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_read_reg2 <= clr_read_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_rstat_reg <= ((end_operation OR do_read_sid) OR do_read);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_rstat_reg2 <= clr_rstat_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_secprot_reg <= (((wire_spstage_cntr_q(1) AND wire_spstage_cntr_q(0)) AND end_operation) OR do_read_sid);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_secprot_reg2 <= clr_secprot_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_write_reg <= ((((((wire_w_lg_w_lg_w586w587w588w(0) OR wire_w_lg_do_write63w(0)) OR wire_w584w(0)) OR do_read_sid) OR do_sec_prot) OR do_read) OR do_fast_read);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_write_reg2 <= clr_write_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN cnt_bfend_reg <= cnt_bfend_wire_in;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN do_wrmemadd_reg <= (wire_wrstage_cntr_q(1) AND wire_wrstage_cntr_q(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, end_operation)
	BEGIN
		IF (end_operation = '1') THEN dvalid_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_dvalid_reg_ena = '1') THEN dvalid_reg <= (end_read_byte AND end_one_cyc_pos);
			END IF;
		END IF;
	END PROCESS;
	wire_dvalid_reg_ena <= wire_w_lg_do_read330w(0);
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN dvalid_reg2 <= dvalid_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN end1_cyc_reg <= end1_cyc_reg_in_wire;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN end1_cyc_reg2 <= end_one_cycle;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN end_op_hdlyreg <= end_operation;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN end_op_reg <= ((((((((((wire_stage_cntr_w_lg_w_q_range89w94w(0) AND ((wire_w_lg_w_lg_w_lg_w_lg_do_read274w275w276w277w(0) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read))) OR (wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range89w92w269w270w(0) AND wire_w_lg_do_polling268w(0))) OR ((((((do_read_rdid AND end_one_cycle) AND wire_stage_cntr_q(1)) AND wire_stage_cntr_q(0)) AND wire_addbyte_cntr_q(2)) AND wire_addbyte_cntr_q(1)) AND wire_addbyte_cntr_q(0))) OR (wire_w_lg_w_lg_start_poll259w260w(0) AND wire_w_lg_st_busy_wire102w(0))) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range89w90w91w257w258w(0)) OR wire_w_lg_w_lg_w_lg_do_write65w66w67w(0)) OR wire_w_lg_w_lg_do_write56w253w(0)) OR wire_w_lg_do_write63w(0)) OR wire_stage_cntr_w252w(0)) OR wire_stage_cntr_w_lg_w247w248w(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN end_opfdly_reg <= end_operation;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN end_pgwrop_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_end_pgwrop_reg_ena = '1') THEN end_pgwrop_reg <= buf_empty;
			END IF;
		END IF;
	END PROCESS;
	wire_end_pgwrop_reg_ena <= ((cnt_bfend_reg AND do_write) AND shift_pgwr_data);
	PROCESS (clkin_wire, clr_endrbyte_reg)
	BEGIN
		IF (clr_endrbyte_reg = '1') THEN end_rbyte_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_end_rbyte_reg_ena = '1') THEN end_rbyte_reg <= wire_w_lg_w_lg_w_lg_do_read330w374w375w(0);
			END IF;
		END IF;
	END PROCESS;
	wire_end_rbyte_reg_ena <= (wire_gen_cntr_w_lg_w_q_range99w100w(0) AND wire_gen_cntr_q(0));
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN end_read_reg <= (((wire_w_lg_rden_wire389w(0) AND wire_w_lg_do_read330w(0)) AND data_valid_wire) AND end_read_byte);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_read_wire)
	BEGIN
		IF (clr_read_wire = '1') THEN fast_read_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_fast_read_reg_ena = '1') THEN fast_read_reg <= fast_read;
			END IF;
		END IF;
	END PROCESS;
	wire_fast_read_reg_ena <= (wire_w_lg_busy_wire2w(0) AND rden_wire);
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN ill_erase_reg <= (illegal_erase_dly_reg OR illegal_erase_b4out_wire);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN ill_write_reg <= (illegal_write_dly_reg OR illegal_write_b4out_wire);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (power_up_reg = '1') THEN illegal_erase_dly_reg <= illegal_erase_b4out_wire;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (power_up_reg = '1') THEN illegal_write_dly_reg <= illegal_write_b4out_wire;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN max_cnt_reg <= wire_cmpr5_aeb;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN maxcnt_shift_reg <= (wire_w_lg_w_lg_reach_max_cnt484w485w(0) AND wire_w_lg_do_write408w(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN maxcnt_shift_reg2 <= maxcnt_shift_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, end_ophdly)
	BEGIN
		IF (end_ophdly = '1') THEN ncs_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_ncs_reg_ena = '1') THEN ncs_reg <= '1';
			END IF;
		END IF;
	END PROCESS;
	wire_ncs_reg_ena <= (wire_stage_cntr_w_lg_w_lg_w_q_range89w90w91w(0) AND end_one_cyc_pos);
	wire_ncs_reg_w_lg_q291w(0) <= NOT ncs_reg;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(0) = '1') THEN pgwrbuf_dataout(0) <= wire_pgwrbuf_dataout_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(1) = '1') THEN pgwrbuf_dataout(1) <= wire_pgwrbuf_dataout_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(2) = '1') THEN pgwrbuf_dataout(2) <= wire_pgwrbuf_dataout_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(3) = '1') THEN pgwrbuf_dataout(3) <= wire_pgwrbuf_dataout_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(4) = '1') THEN pgwrbuf_dataout(4) <= wire_pgwrbuf_dataout_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(5) = '1') THEN pgwrbuf_dataout(5) <= wire_pgwrbuf_dataout_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(6) = '1') THEN pgwrbuf_dataout(6) <= wire_pgwrbuf_dataout_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(7) = '1') THEN pgwrbuf_dataout(7) <= wire_pgwrbuf_dataout_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_pgwrbuf_dataout_d <= ( wire_w_lg_w_lg_read_bufdly442w443w & wire_w_lg_read_bufdly447w);
	loop34 : FOR i IN 0 TO 7 GENERATE
		wire_pgwrbuf_dataout_ena(i) <= wire_w_lg_read_bufdly437w(0);
	END GENERATE loop34;
	wire_pgwrbuf_dataout_w_q_range438w <= pgwrbuf_dataout(6 DOWNTO 0);
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN power_up_reg <= (busy_wire OR busy_delay_reg);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (rdid_load = '1') THEN rdid_out_reg <= ( read_dout_reg(7 DOWNTO 0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN read_bufdly_reg <= read_buf;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(0) = '1') THEN read_data_reg(0) <= wire_read_data_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(1) = '1') THEN read_data_reg(1) <= wire_read_data_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(2) = '1') THEN read_data_reg(2) <= wire_read_data_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(3) = '1') THEN read_data_reg(3) <= wire_read_data_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(4) = '1') THEN read_data_reg(4) <= wire_read_data_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(5) = '1') THEN read_data_reg(5) <= wire_read_data_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(6) = '1') THEN read_data_reg(6) <= wire_read_data_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(7) = '1') THEN read_data_reg(7) <= wire_read_data_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_read_data_reg_d <= ( read_data_reg_in_wire(7 DOWNTO 0));
	loop35 : FOR i IN 0 TO 7 GENERATE
		wire_read_data_reg_ena(i) <= wire_w377w(0);
	END GENERATE loop35;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(0) = '1') THEN read_dout_reg(0) <= wire_read_dout_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(1) = '1') THEN read_dout_reg(1) <= wire_read_dout_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(2) = '1') THEN read_dout_reg(2) <= wire_read_dout_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(3) = '1') THEN read_dout_reg(3) <= wire_read_dout_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(4) = '1') THEN read_dout_reg(4) <= wire_read_dout_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(5) = '1') THEN read_dout_reg(5) <= wire_read_dout_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(6) = '1') THEN read_dout_reg(6) <= wire_read_dout_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(7) = '1') THEN read_dout_reg(7) <= wire_read_dout_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_read_dout_reg_d <= ( read_dout_reg(6 DOWNTO 0) & wire_w_lg_data0out_wire346w);
	loop36 : FOR i IN 0 TO 7 GENERATE
		wire_read_dout_reg_ena(i) <= wire_w_lg_w_lg_stage4_wire343w344w(0);
	END GENERATE loop36;
	PROCESS (clkin_wire, clr_rdid_wire)
	BEGIN
		IF (clr_rdid_wire = '1') THEN read_rdid_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (busy_wire = '0') THEN read_rdid_reg <= read_rdid;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN read_status_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (busy_wire = '0') THEN read_status_reg <= read_status;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN sec_erase_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_sec_erase_reg_ena = '1') THEN sec_erase_reg <= sector_erase;
			END IF;
		END IF;
	END PROCESS;
	wire_sec_erase_reg_ena <= (wire_w_lg_busy_wire2w(0) AND wren_wire);
	PROCESS (clkin_wire, clr_secprot_wire)
	BEGIN
		IF (clr_secprot_wire = '1') THEN sec_prot_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_sec_prot_reg_ena = '1') THEN sec_prot_reg <= sector_protect;
			END IF;
		END IF;
	END PROCESS;
	wire_sec_prot_reg_ena <= (wire_w_lg_busy_wire2w(0) AND wren_wire);
	PROCESS (clkin_wire, end_ophdly)
	BEGIN
		IF (end_ophdly = '1') THEN shftpgwr_data_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN shftpgwr_data_reg <= ((wire_stage_cntr_w_lg_w_q_range89w94w(0) AND wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_q(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN shift_op_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range89w90w91w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_secprot_wire)
	BEGIN
		IF (clr_secprot_wire = '1') THEN sprot_rstat_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN sprot_rstat_reg <= (wire_w_lg_do_sec_prot621w(0) AND wire_spstage_cntr_q(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN stage2_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range89w90w91w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN stage3_dly_reg <= wire_stage_cntr_w_lg_w_q_range89w92w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN stage3_reg <= wire_stage_cntr_w_lg_w_q_range89w92w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN stage4_reg <= wire_stage_cntr_w_lg_w_q_range89w94w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_secprot_wire)
	BEGIN
		IF (clr_secprot_wire = '1') THEN start_sppoll_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_start_sppoll_reg_ena = '1') THEN start_sppoll_reg <= wire_stage_cntr_w_lg_w_q_range89w92w(0);
			END IF;
		END IF;
	END PROCESS;
	wire_start_sppoll_reg_ena <= ((do_sprot_rstat AND do_polling) AND end_one_cycle);
	PROCESS (clkin_wire, clr_secprot_wire)
	BEGIN
		IF (clr_secprot_wire = '1') THEN start_sppoll_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN start_sppoll_reg2 <= start_sppoll_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN start_wrpoll_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_start_wrpoll_reg_ena = '1') THEN start_wrpoll_reg <= wire_stage_cntr_w_lg_w_q_range89w92w(0);
			END IF;
		END IF;
	END PROCESS;
	wire_start_wrpoll_reg_ena <= ((do_write_rstat AND do_polling) AND end_one_cycle);
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN start_wrpoll_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN start_wrpoll_reg2 <= start_wrpoll_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(0) = '1') THEN statreg_int(0) <= wire_statreg_int_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(1) = '1') THEN statreg_int(1) <= wire_statreg_int_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(2) = '1') THEN statreg_int(2) <= wire_statreg_int_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(3) = '1') THEN statreg_int(3) <= wire_statreg_int_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(4) = '1') THEN statreg_int(4) <= wire_statreg_int_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(5) = '1') THEN statreg_int(5) <= wire_statreg_int_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(6) = '1') THEN statreg_int(6) <= wire_statreg_int_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(7) = '1') THEN statreg_int(7) <= wire_statreg_int_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_statreg_int_d <= ( read_dout_reg(7 DOWNTO 0));
	loop37 : FOR i IN 0 TO 7 GENERATE
		wire_statreg_int_ena(i) <= wire_w_lg_w_lg_end_operation422w423w(0);
	END GENERATE loop37;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(0) = '1') THEN statreg_out(0) <= wire_statreg_out_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(1) = '1') THEN statreg_out(1) <= wire_statreg_out_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(2) = '1') THEN statreg_out(2) <= wire_statreg_out_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(3) = '1') THEN statreg_out(3) <= wire_statreg_out_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(4) = '1') THEN statreg_out(4) <= wire_statreg_out_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(5) = '1') THEN statreg_out(5) <= wire_statreg_out_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(6) = '1') THEN statreg_out(6) <= wire_statreg_out_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(7) = '1') THEN statreg_out(7) <= wire_statreg_out_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_statreg_out_d <= ( read_dout_reg(7 DOWNTO 0));
	loop38 : FOR i IN 0 TO 7 GENERATE
		wire_statreg_out_ena(i) <= wire_w_lg_w413w414w(0);
	END GENERATE loop38;
	PROCESS (clkin_wire, end_opfdly)
	BEGIN
		IF (end_opfdly = '1') THEN streg_datain_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_streg_datain_reg_ena = '1') THEN streg_datain_reg <= wrstat_dreg(7);
			END IF;
		END IF;
	END PROCESS;
	wire_streg_datain_reg_ena <= (wire_w_lg_do_sec_prot600w(0) AND wire_spstage_cntr_q(0));
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN write_prot_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_write_prot_reg_ena = '1') THEN write_prot_reg <= ((wire_w_lg_do_write65w(0) AND (((((wire_addr_reg_w_lg_w_lg_w535w536w537w(0) OR (wire_addr_reg_w531w(0) AND wire_w_lg_bp0_wire516w(0))) OR wire_addr_reg_w527w(0)) OR ((wire_addr_reg_w_lg_w_lg_w_q_range512w518w519w(0) AND wire_w_lg_bp1_wire511w(0)) AND wire_w_lg_bp0_wire516w(0))) OR wire_addr_reg_w_lg_w_lg_w_lg_w_q_range512w513w514w515w(0)) OR (bp2_wire AND bp1_wire))) OR be_write_prot);
			END IF;
		END IF;
	END PROCESS;
	wire_write_prot_reg_ena <= (((wire_w_lg_w_lg_do_sec_erase501w502w(0) AND (NOT wire_wrstage_cntr_q(1))) AND wire_wrstage_cntr_q(0)) AND end_ophdly);
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN write_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_write_reg_ena = '1') THEN write_reg <= write;
			END IF;
		END IF;
	END PROCESS;
	wire_write_reg_ena <= (wire_w_lg_busy_wire2w(0) AND wren_wire);
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN write_rstat_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN write_rstat_reg <= (wire_w_lg_w_lg_w_lg_do_write65w66w499w(0) AND (((NOT wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_w_lg_w_q_range492w493w(0)) OR wire_wrstage_cntr_w_lg_w_q_range494w495w(0)));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_secprot_wire)
	BEGIN
		IF (clr_secprot_wire = '1') THEN wrstat_dreg(0) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_wrstat_dreg_ena(0) = '1') THEN wrstat_dreg(0) <= wire_wrstat_dreg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_secprot_wire)
	BEGIN
		IF (clr_secprot_wire = '1') THEN wrstat_dreg(1) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_wrstat_dreg_ena(1) = '1') THEN wrstat_dreg(1) <= wire_wrstat_dreg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_secprot_wire)
	BEGIN
		IF (clr_secprot_wire = '1') THEN wrstat_dreg(2) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_wrstat_dreg_ena(2) = '1') THEN wrstat_dreg(2) <= wire_wrstat_dreg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_secprot_wire)
	BEGIN
		IF (clr_secprot_wire = '1') THEN wrstat_dreg(3) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_wrstat_dreg_ena(3) = '1') THEN wrstat_dreg(3) <= wire_wrstat_dreg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_secprot_wire)
	BEGIN
		IF (clr_secprot_wire = '1') THEN wrstat_dreg(4) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_wrstat_dreg_ena(4) = '1') THEN wrstat_dreg(4) <= wire_wrstat_dreg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_secprot_wire)
	BEGIN
		IF (clr_secprot_wire = '1') THEN wrstat_dreg(5) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_wrstat_dreg_ena(5) = '1') THEN wrstat_dreg(5) <= wire_wrstat_dreg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_secprot_wire)
	BEGIN
		IF (clr_secprot_wire = '1') THEN wrstat_dreg(6) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_wrstat_dreg_ena(6) = '1') THEN wrstat_dreg(6) <= wire_wrstat_dreg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_secprot_wire)
	BEGIN
		IF (clr_secprot_wire = '1') THEN wrstat_dreg(7) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_wrstat_dreg_ena(7) = '1') THEN wrstat_dreg(7) <= wire_wrstat_dreg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_wrstat_dreg_d <= ( wire_w_lg_w_lg_not_busy605w606w & wire_w_lg_not_busy610w);
	loop39 : FOR i IN 0 TO 7 GENERATE
		wire_wrstat_dreg_ena(i) <= wire_w_lg_w_lg_wren_wire615w616w(0);
	END GENERATE loop39;
	wire_wrstat_dreg_w_q_range602w <= wrstat_dreg(6 DOWNTO 0);
	wire_cmpr5_dataa <= ( page_size_wire(8 DOWNTO 0));
	wire_cmpr5_datab <= ( wire_pgwr_data_cntr_q(8 DOWNTO 0));
	cmpr5 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aeb => wire_cmpr5_aeb,
		dataa => wire_cmpr5_dataa,
		datab => wire_cmpr5_datab
	  );
	wire_cmpr6_dataa <= ( wire_pgwr_data_cntr_q(8 DOWNTO 0));
	wire_cmpr6_datab <= ( wire_pgwr_read_cntr_q(8 DOWNTO 0));
	cmpr6 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aeb => wire_cmpr6_aeb,
		dataa => wire_cmpr6_dataa,
		datab => wire_cmpr6_datab
	  );
	wire_pgwr_data_cntr_clk_en <= wire_w_lg_w_lg_w_lg_shift_bytes_wire434w450w451w(0);
	wire_w_lg_w_lg_w_lg_shift_bytes_wire434w450w451w(0) <= ((shift_bytes_wire AND wren_wire) AND wire_w_lg_reach_max_cnt449w(0)) AND wire_w_lg_do_write408w(0);
	wire_pgwr_data_cntr_w_q_range455w(0) <= wire_pgwr_data_cntr_q(1);
	wire_pgwr_data_cntr_w_q_range458w(0) <= wire_pgwr_data_cntr_q(2);
	wire_pgwr_data_cntr_w_q_range461w(0) <= wire_pgwr_data_cntr_q(3);
	wire_pgwr_data_cntr_w_q_range464w(0) <= wire_pgwr_data_cntr_q(4);
	wire_pgwr_data_cntr_w_q_range467w(0) <= wire_pgwr_data_cntr_q(5);
	wire_pgwr_data_cntr_w_q_range470w(0) <= wire_pgwr_data_cntr_q(6);
	wire_pgwr_data_cntr_w_q_range473w(0) <= wire_pgwr_data_cntr_q(7);
	wire_pgwr_data_cntr_w_q_range476w(0) <= wire_pgwr_data_cntr_q(8);
	pgwr_data_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 9
	  )
	  PORT MAP ( 
		aclr => clr_write_wire,
		clk_en => wire_pgwr_data_cntr_clk_en,
		clock => clkin_wire,
		q => wire_pgwr_data_cntr_q
	  );
	pgwr_read_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 9
	  )
	  PORT MAP ( 
		aclr => clr_write_wire,
		clk_en => read_buf,
		clock => clkin_wire,
		q => wire_pgwr_read_cntr_q
	  );
	wire_mux211_dataout <= end1_cyc_dlyncs_in_wire WHEN (((do_write OR do_sec_prot) OR do_sec_erase) OR do_bulk_erase) = '1'  ELSE end1_cyc_normal_in_wire;
	wire_mux212_dataout <= end_add_cycle_mux_datab_wire WHEN do_fast_read = '1'  ELSE wire_addbyte_cntr_w_lg_w_q_range137w142w(0);
	wire_scfifo4_data <= ( datain(7 DOWNTO 0));
	wire_scfifo4_rdreq <= wire_w_lg_read_buf436w(0);
	wire_w_lg_read_buf436w(0) <= read_buf OR dummy_read_buf;
	wire_scfifo4_wrreq <= wire_w_lg_w_lg_shift_bytes_wire434w435w(0);
	wire_w_lg_w_lg_shift_bytes_wire434w435w(0) <= (shift_bytes_wire AND wren_wire) AND wire_w_lg_do_write408w(0);
	wire_scfifo4_w_q_range441w <= wire_scfifo4_q(7 DOWNTO 1);
	wire_scfifo4_w_q_range446w(0) <= wire_scfifo4_q(0);
	scfifo4 :  scfifo
	  GENERIC MAP (
		LPM_NUMWORDS => 258,
		LPM_WIDTH => 8,
		LPM_WIDTHU => 9,
		USE_EAB => "ON"
	  )
	  PORT MAP ( 
		aclr => clr_write_wire,
		clock => clkin_wire,
		data => wire_scfifo4_data,
		q => wire_scfifo4_q,
		rdreq => wire_scfifo4_rdreq,
		wrreq => wire_scfifo4_wrreq
	  );

 END RTL; --z126_01_pasmi_sim_m25p32_altasmi_parallel_l2q2
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY z126_01_pasmi_sim_m25p32 IS
	PORT
	(
		addr		: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
		bulk_erase		: IN STD_LOGIC ;
		clkin		: IN STD_LOGIC ;
		datain		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		fast_read		: IN STD_LOGIC ;
		rden		: IN STD_LOGIC ;
		read_rdid		: IN STD_LOGIC ;
		read_status		: IN STD_LOGIC ;
		sector_erase		: IN STD_LOGIC ;
		sector_protect		: IN STD_LOGIC ;
		shift_bytes		: IN STD_LOGIC ;
		wren		: IN STD_LOGIC ;
		write		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		data_valid		: OUT STD_LOGIC ;
		dataout		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		illegal_erase		: OUT STD_LOGIC ;
		illegal_write		: OUT STD_LOGIC ;
		rdid_out		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		status_out		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END z126_01_pasmi_sim_m25p32;


ARCHITECTURE RTL OF z126_01_pasmi_sim_m25p32 IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "ALTASMI_PARALLEL";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "data_width=STANDARD;epcs_type=EPCS16;intended_device_family=Cyclone III;lpm_hint=UNUSED;lpm_type=altasmi_parallel;page_size=256;port_bulk_erase=PORT_USED;port_en4b_addr=PORT_UNUSED;port_fast_read=PORT_USED;port_illegal_erase=PORT_USED;port_illegal_write=PORT_USED;port_rdid_out=PORT_USED;port_read_address=PORT_UNUSED;port_read_rdid=PORT_USED;port_read_sid=PORT_UNUSED;port_read_status=PORT_USED;port_sector_erase=PORT_USED;port_sector_protect=PORT_USED;port_shift_bytes=PORT_USED;port_wren=PORT_USED;port_write=PORT_USED;use_eab=ON;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC ;
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC ;



	COMPONENT z126_01_pasmi_sim_m25p32_altasmi_parallel_l2q2
	PORT (
			sector_protect	: IN STD_LOGIC ;
			bulk_erase	: IN STD_LOGIC ;
			clkin	: IN STD_LOGIC ;
			data_valid	: OUT STD_LOGIC ;
			datain	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			fast_read	: IN STD_LOGIC ;
			illegal_erase	: OUT STD_LOGIC ;
			rden	: IN STD_LOGIC ;
			dataout	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			rdid_out	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			read_rdid	: IN STD_LOGIC ;
			addr	: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
			busy	: OUT STD_LOGIC ;
			read_status	: IN STD_LOGIC ;
			sector_erase	: IN STD_LOGIC ;
			status_out	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			write	: IN STD_LOGIC ;
			illegal_write	: OUT STD_LOGIC ;
			shift_bytes	: IN STD_LOGIC ;
			wren	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	data_valid    <= sub_wire0;
	illegal_erase    <= sub_wire1;
	dataout    <= sub_wire2(7 DOWNTO 0);
	rdid_out    <= sub_wire3(7 DOWNTO 0);
	busy    <= sub_wire4;
	status_out    <= sub_wire5(7 DOWNTO 0);
	illegal_write    <= sub_wire6;

	z126_01_pasmi_sim_m25p32_altasmi_parallel_l2q2_component : z126_01_pasmi_sim_m25p32_altasmi_parallel_l2q2
	PORT MAP (
		sector_protect => sector_protect,
		bulk_erase => bulk_erase,
		clkin => clkin,
		datain => datain,
		fast_read => fast_read,
		rden => rden,
		read_rdid => read_rdid,
		addr => addr,
		read_status => read_status,
		sector_erase => sector_erase,
		write => write,
		shift_bytes => shift_bytes,
		wren => wren,
		data_valid => sub_wire0,
		illegal_erase => sub_wire1,
		dataout => sub_wire2,
		rdid_out => sub_wire3,
		busy => sub_wire4,
		status_out => sub_wire5,
		illegal_write => sub_wire6
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
-- Retrieval info: CONSTANT: DATA_WIDTH STRING "STANDARD"
-- Retrieval info: CONSTANT: EPCS_TYPE STRING "EPCS16"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altasmi_parallel"
-- Retrieval info: CONSTANT: PAGE_SIZE NUMERIC "256"
-- Retrieval info: CONSTANT: PORT_BULK_ERASE STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_EN4B_ADDR STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_FAST_READ STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_ILLEGAL_ERASE STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_ILLEGAL_WRITE STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_RDID_OUT STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_READ_ADDRESS STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_RDID STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_READ_SID STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_STATUS STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_SECTOR_ERASE STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_SECTOR_PROTECT STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_SHIFT_BYTES STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_WREN STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_WRITE STRING "PORT_USED"
-- Retrieval info: CONSTANT: USE_EAB STRING "ON"
-- Retrieval info: USED_PORT: addr 0 0 24 0 INPUT NODEFVAL "addr[23..0]"
-- Retrieval info: CONNECT: @addr 0 0 24 0 addr 0 0 24 0
-- Retrieval info: USED_PORT: bulk_erase 0 0 0 0 INPUT NODEFVAL "bulk_erase"
-- Retrieval info: CONNECT: @bulk_erase 0 0 0 0 bulk_erase 0 0 0 0
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: USED_PORT: clkin 0 0 0 0 INPUT NODEFVAL "clkin"
-- Retrieval info: CONNECT: @clkin 0 0 0 0 clkin 0 0 0 0
-- Retrieval info: USED_PORT: data_valid 0 0 0 0 OUTPUT NODEFVAL "data_valid"
-- Retrieval info: CONNECT: data_valid 0 0 0 0 @data_valid 0 0 0 0
-- Retrieval info: USED_PORT: datain 0 0 8 0 INPUT NODEFVAL "datain[7..0]"
-- Retrieval info: CONNECT: @datain 0 0 8 0 datain 0 0 8 0
-- Retrieval info: USED_PORT: dataout 0 0 8 0 OUTPUT NODEFVAL "dataout[7..0]"
-- Retrieval info: CONNECT: dataout 0 0 8 0 @dataout 0 0 8 0
-- Retrieval info: USED_PORT: fast_read 0 0 0 0 INPUT NODEFVAL "fast_read"
-- Retrieval info: CONNECT: @fast_read 0 0 0 0 fast_read 0 0 0 0
-- Retrieval info: USED_PORT: illegal_erase 0 0 0 0 OUTPUT NODEFVAL "illegal_erase"
-- Retrieval info: CONNECT: illegal_erase 0 0 0 0 @illegal_erase 0 0 0 0
-- Retrieval info: USED_PORT: illegal_write 0 0 0 0 OUTPUT NODEFVAL "illegal_write"
-- Retrieval info: CONNECT: illegal_write 0 0 0 0 @illegal_write 0 0 0 0
-- Retrieval info: USED_PORT: rden 0 0 0 0 INPUT NODEFVAL "rden"
-- Retrieval info: CONNECT: @rden 0 0 0 0 rden 0 0 0 0
-- Retrieval info: USED_PORT: rdid_out 0 0 8 0 OUTPUT NODEFVAL "rdid_out[7..0]"
-- Retrieval info: CONNECT: rdid_out 0 0 8 0 @rdid_out 0 0 8 0
-- Retrieval info: USED_PORT: read_rdid 0 0 0 0 INPUT NODEFVAL "read_rdid"
-- Retrieval info: CONNECT: @read_rdid 0 0 0 0 read_rdid 0 0 0 0
-- Retrieval info: USED_PORT: read_status 0 0 0 0 INPUT NODEFVAL "read_status"
-- Retrieval info: CONNECT: @read_status 0 0 0 0 read_status 0 0 0 0
-- Retrieval info: USED_PORT: sector_erase 0 0 0 0 INPUT NODEFVAL "sector_erase"
-- Retrieval info: CONNECT: @sector_erase 0 0 0 0 sector_erase 0 0 0 0
-- Retrieval info: USED_PORT: sector_protect 0 0 0 0 INPUT NODEFVAL "sector_protect"
-- Retrieval info: CONNECT: @sector_protect 0 0 0 0 sector_protect 0 0 0 0
-- Retrieval info: USED_PORT: shift_bytes 0 0 0 0 INPUT NODEFVAL "shift_bytes"
-- Retrieval info: CONNECT: @shift_bytes 0 0 0 0 shift_bytes 0 0 0 0
-- Retrieval info: USED_PORT: status_out 0 0 8 0 OUTPUT NODEFVAL "status_out[7..0]"
-- Retrieval info: CONNECT: status_out 0 0 8 0 @status_out 0 0 8 0
-- Retrieval info: USED_PORT: wren 0 0 0 0 INPUT NODEFVAL "wren"
-- Retrieval info: CONNECT: @wren 0 0 0 0 wren 0 0 0 0
-- Retrieval info: USED_PORT: write 0 0 0 0 INPUT NODEFVAL "write"
-- Retrieval info: CONNECT: @write 0 0 0 0 write 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL z126_01_pasmi_sim_m25p32_2.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL z126_01_pasmi_sim_m25p32_2.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL z126_01_pasmi_sim_m25p32_2.bsf FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL z126_01_pasmi_sim_m25p32_2_inst.vhd FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL z126_01_pasmi_sim_m25p32_2.inc FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL z126_01_pasmi_sim_m25p32_2.cmp FALSE TRUE

